module patch (w98, n29, n31, n33, n36);
input n29, n31, n33, n36;
output w98;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98;
not(w0, n31);
not(w1, n33);
or (w2, n29, n36);
or (w3, w0, n36);
or (w4, w1, n36);
and (w5, w3, w4);
and (w6, w5, w2);
and (w7, w2, w3);
and (w8, w7, w6);
and (w9, w6, w2);
and (w10, w8, w9);
and (w11, w10, w9);
and (w12, w11, w2);
and (w13, w7, w12);
and (w14, w13, w9);
and (w15, w14, w9);
and (w16, w15, w2);
and (w17, w4, w3);
and (w18, w17, w2);
and (w19, w18, w16);
and (w20, w19, w9);
and (w21, w20, w2);
and (w22, w21, w20);
and (w23, w22, w20);
and (w24, w23, w18);
and (w25, w24, w20);
and (w26, w2, w20);
and (w27, w26, w20);
and (w28, w27, w20);
and (w29, w28, w20);
and (w30, w29, w25);
and (w31, w30, w20);
and (w32, w31, w18);
and (w33, w32, w20);
and (w34, w33, w18);
and (w35, w34, w33);
and (w36, w35, w8);
and (w37, w36, w35);
and (w38, w37, w33);
and (w39, w38, w33);
and (w40, w39, w33);
and (w41, w40, w33);
and (w42, w41, w20);
and (w43, w42, w33);
and (w44, w43, w33);
and (w45, w44, w33);
and (w46, w45, w20);
and (w47, w46, w33);
and (w48, w47, w2);
and (w49, w48, w2);
and (w50, w49, w2);
and (w51, w33, w7);
and (w52, w51, w35);
and (w53, w52, w33);
and (w54, w53, w33);
and (w55, w54, w33);
and (w56, w55, w35);
and (w57, w56, w33);
and (w58, w57, w33);
and (w59, w58, w20);
and (w60, w59, w33);
and (w61, w60, w33);
and (w62, w61, w20);
and (w63, w55, w35);
and (w64, w63, w33);
and (w65, w64, w33);
and (w66, w65, w33);
and (w67, w66, w20);
and (w68, w67, w33);
and (w69, w68, w20);
and (w70, w69, w62);
and (w71, w33, w50);
and (w72, w71, w50);
and (w73, w72, w2);
and (w74, w33, w50);
and (w75, w74, w50);
and (w76, w75, w20);
and (w77, w76, w20);
and (w78, w77, w73);
and (w79, w33, w50);
and (w80, w79, w50);
and (w81, w80, w78);
and (w82, w81, w20);
and (w83, w82, w20);
and (w84, w83, w73);
and (w85, w70, w84);
and (w86, w85, w33);
and (w87, w86, w33);
and (w88, w87, w2);
and (w89, w88, w2);
and (w90, w89, w20);
and (w91, w89, w20);
and (w92, w2, w85);
and (w93, w92, w90);
and (w94, w93, w91);
and (w95, w94, w33);
and (w96, w94, w33);
and (w97, w95, w85);
and (w98, w97, w96);
endmodule