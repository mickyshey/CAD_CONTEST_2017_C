module patch (w23, a, b, c);
input a, b, c;
output w23;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23;
or (w0, !b, !c);
and (w1, a, !a);
or (w2, w1, c);
and (w3, w2, w0);
or (w4, w3, !b);
and (w5, w4, b);
or (w6, w5, !c);
or (w7, w6, !c);
or (w8, w7, !a);
or (w9, w8, b);
and (w10, !b, w9);
and (w11, !b, w9);
or (w12, w10, w5);
and (w13, c, w9);
or (w14, w13, w11);
or (w15, w14, w12);
or (w16, a, w15);
and (w17, w16, w9);
and (w18, w16, w9);
and (w19, w16, w9);
and (w20, w17, w19);
and (w21, w18, w9);
and (w22, w21, w20);
and (w23, w22, w18);
endmodule