module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 ;
output g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , 
     n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , 
     n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , 
     n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , 
     n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , 
     n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , 
     n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , 
     n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , 
     n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
     n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
     n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
     n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , 
     n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , 
     n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , 
     n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , 
     n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , 
     n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , 
     n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , 
     n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , 
     n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , 
     n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , 
     n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , 
     n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , 
     n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
     n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
     n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
     n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
     n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
     n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
     n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
     n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
     n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
     n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
     n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
     n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
     n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
     n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
     n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
     n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
     n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
     n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , 
     n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
     n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
     n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
     n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
     n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
     n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
     n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
     n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
     n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
     n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
     n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
     n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
     n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
     n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
     n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
     n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
     n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
     n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
     n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
     n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , 
     n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , 
     n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , 
     n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , 
     n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , 
     n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , 
     n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , 
     n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , 
     n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , 
     n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , 
     n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , 
     n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
     n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
     n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
     n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , 
     n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , 
     n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
     n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
     n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
     n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
     n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
     n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
     n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
     n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
     n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
     n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
     n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
     n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
     n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
     n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
     n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
     n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
     n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
     n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
     n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
     n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
     n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
     n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
     n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
     n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
     n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
     n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
     n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
     n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
     n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , 
     n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
     n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
     n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
     n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
     n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
     n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
     n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
     n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
     n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
     n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
     n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
     n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
     n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
     n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
     n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
     n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
     n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
     n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
     n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
     n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , 
     n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , 
     n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
     n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
     n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , 
     n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , 
     n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , 
     n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
     n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
     n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
     n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
     n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
     n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
     n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
     n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
     n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
     n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
     n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
     n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
     n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
     n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , 
     n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , 
     n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , 
     n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , 
     n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , 
     n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , 
     n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , 
     n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , 
     n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
     n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
     n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
     n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
     n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
     n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
     n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , 
     n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , 
     n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , 
     n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , 
     n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , 
     n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
     n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , 
     n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , 
     n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , 
     n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , 
     n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , 
     n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , 
     n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , 
     n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , 
     n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
     n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
     n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
     n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
     n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , 
     n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , 
     n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , 
     n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , 
     n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
     n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
     n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
     n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
     n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , 
     n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
     n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
     n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
     n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
     n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , 
     n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
     n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
     n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
     n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
     n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , 
     n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , 
     n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , 
     n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , 
     n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , 
     n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
     n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , 
     n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , 
     n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , 
     n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
     n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
     n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
     n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
     n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
     n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
     n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
     n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
     n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , 
     n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
     n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
     n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
     n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , 
     n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , 
     n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , 
     n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , 
     n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , 
     n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , 
     n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , 
     n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , 
     n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , 
     n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , 
     n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , 
     n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , 
     n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , 
     n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , 
     n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
     n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , 
     n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , 
     n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , 
     n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
     n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
     n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
     n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
     n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
     n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , 
     n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , 
     n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , 
     n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , 
     n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
     n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
     n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
     n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
     n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
     n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
     n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
     n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
     n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
     n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
     n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
     n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
     n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
     n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
     n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , 
     n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , 
     n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , 
     n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , 
     n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , 
     n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , 
     n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , 
     n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , 
     n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , 
     n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , 
     n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , 
     n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , 
     n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , 
     n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , 
     n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , 
     n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , 
     n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , 
     n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , 
     n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , 
     n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , 
     n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , 
     n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , 
     n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , 
     n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , 
     n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , 
     n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
     n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , 
     n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
     n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
     n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
     n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
     n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
     n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
     n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
     n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
     n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
     n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
     n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
     n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
     n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
     n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
     n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
     n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , 
     n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , 
     n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , 
     n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , 
     n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , 
     n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , 
     n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , 
     n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 ;
wire t_0 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( g46 , n47 );
buf ( g47 , n48 );
buf ( g48 , n49 );
buf ( g49 , n50 );
buf ( g50 , n51 );
buf ( g51 , n52 );
buf ( g52 , n53 );
buf ( g53 , n54 );
buf ( g54 , n55 );
buf ( g55 , n56 );
buf ( g56 , n57 );
buf ( g57 , n58 );
buf ( g58 , n59 );
buf ( g59 , n60 );
buf ( g60 , n61 );
buf ( g61 , n62 );
buf ( g62 , n63 );
buf ( g63 , n64 );
buf ( g64 , n65 );
buf ( g65 , n66 );
buf ( g66 , n67 );
buf ( g67 , n68 );
buf ( g68 , n69 );
buf ( g69 , n70 );
buf ( g70 , n71 );
buf ( g71 , n72 );
buf ( g72 , n73 );
buf ( n47 , n4279 );
buf ( n48 , n7295 );
buf ( n49 , n12680 );
buf ( n50 , n9232 );
buf ( n51 , n11383 );
buf ( n52 , n13778 );
buf ( n53 , n13646 );
buf ( n54 , n12982 );
buf ( n55 , n13015 );
buf ( n56 , n12999 );
buf ( n57 , n13301 );
buf ( n58 , n13354 );
buf ( n59 , n13777 );
buf ( n60 , n13601 );
buf ( n61 , n13453 );
buf ( n62 , n13420 );
buf ( n63 , n13730 );
buf ( n64 , n13231 );
buf ( n65 , n13676 );
buf ( n66 , n13507 );
buf ( n67 , n13763 );
buf ( n68 , n13671 );
buf ( n69 , n13770 );
buf ( n70 , n4225 );
buf ( n71 , n13754 );
buf ( n72 , n13696 );
buf ( n73 , n13775 );
not ( n76 , n13 );
not ( n77 , n2 );
nand ( n78 , n11 , n77 );
nor ( n79 , n12 , n78 );
and ( n80 , n76 , n79 );
not ( n81 , n80 );
nor ( n82 , n20 , n81 );
nor ( n83 , n40 , n41 );
not ( n84 , n83 );
not ( n85 , n84 );
not ( n86 , n85 );
not ( n87 , n86 );
not ( n88 , n87 );
not ( n89 , n88 );
buf ( n90 , n89 );
not ( n91 , n19 );
not ( n92 , n15 );
nand ( n93 , n16 , n17 );
or ( n94 , n92 , n93 );
not ( n95 , n94 );
and ( n96 , n14 , n95 );
and ( n97 , n91 , n96 );
not ( n98 , n97 );
nor ( n99 , n90 , n98 );
nand ( n100 , n22 , n23 );
buf ( n101 , n100 );
not ( n102 , n101 );
not ( n103 , n102 );
not ( n104 , n23 );
nand ( n105 , n104 , n21 , n22 );
and ( n106 , n103 , n105 );
not ( n107 , n22 );
nor ( n108 , n23 , n31 );
not ( n109 , n108 );
not ( n110 , n109 );
nand ( n111 , n107 , n110 );
not ( n112 , n111 );
not ( n113 , n24 );
and ( n114 , n21 , n113 );
not ( n115 , n24 );
not ( n116 , n26 );
nor ( n117 , n116 , n25 );
not ( n118 , n117 );
not ( n119 , n118 );
not ( n120 , n29 );
not ( n121 , n27 );
nor ( n122 , n121 , n28 );
and ( n123 , n120 , n122 );
not ( n124 , n120 );
not ( n125 , n27 );
and ( n126 , n125 , n30 );
nor ( n127 , n126 , n28 );
and ( n128 , n124 , n127 );
nor ( n129 , n123 , n128 );
not ( n130 , n129 );
or ( n131 , n119 , n130 );
not ( n132 , n27 );
nor ( n133 , n132 , n28 );
not ( n134 , n133 );
nand ( n135 , n134 , n117 );
nand ( n136 , n131 , n135 );
nand ( n137 , n115 , n136 );
nand ( n138 , n112 , n114 , n137 );
nand ( n139 , n106 , n138 );
not ( n140 , n139 );
not ( n141 , n21 );
nor ( n142 , n141 , n137 );
buf ( n143 , n142 );
not ( n144 , n143 );
buf ( n145 , n144 );
not ( n146 , n145 );
not ( n147 , n146 );
not ( n148 , n110 );
not ( n149 , n148 );
not ( n150 , n149 );
not ( n151 , n150 );
not ( n152 , n151 );
not ( n153 , n152 );
not ( n154 , n153 );
not ( n155 , n35 );
not ( n156 , n32 );
nand ( n157 , n25 , n33 );
not ( n158 , n157 );
not ( n159 , n158 );
not ( n160 , n159 );
not ( n161 , n160 );
not ( n162 , n161 );
not ( n163 , n162 );
not ( n164 , n127 );
not ( n165 , n34 );
buf ( n166 , n29 );
and ( n167 , n164 , n165 , n166 );
not ( n168 , n167 );
nor ( n169 , n29 , n30 );
not ( n170 , n169 );
not ( n171 , n28 );
not ( n172 , n171 );
or ( n173 , n170 , n172 );
not ( n174 , n34 );
nand ( n175 , n173 , n174 );
not ( n176 , n34 );
nand ( n177 , n176 , n36 );
nand ( n178 , n175 , n177 );
not ( n179 , n178 );
not ( n180 , n179 );
buf ( n181 , n129 );
nand ( n182 , n180 , n181 );
nand ( n183 , n168 , n182 );
not ( n184 , n183 );
not ( n185 , n129 );
not ( n186 , n185 );
nand ( n187 , n186 , n34 );
not ( n188 , n187 );
nor ( n189 , n30 , n36 );
not ( n190 , n29 );
not ( n191 , n190 );
not ( n192 , n191 );
and ( n193 , n178 , n189 , n192 );
nor ( n194 , n188 , n193 );
nand ( n195 , n184 , n194 );
not ( n196 , n195 );
or ( n197 , n163 , n196 );
not ( n198 , n33 );
and ( n199 , n198 , n25 );
not ( n200 , n199 );
not ( n201 , n200 );
not ( n202 , n201 );
not ( n203 , n202 );
and ( n204 , n34 , n181 );
not ( n205 , n34 );
buf ( n206 , n164 );
and ( n207 , n205 , n206 );
nor ( n208 , n204 , n207 );
not ( n209 , n208 );
nand ( n210 , n203 , n209 );
nand ( n211 , n197 , n210 );
nand ( n212 , n156 , n211 );
not ( n213 , n33 );
nor ( n214 , n26 , n32 );
nand ( n215 , n37 , n213 , n214 );
not ( n216 , n215 );
not ( n217 , n209 );
not ( n218 , n217 );
nand ( n219 , n216 , n218 );
nor ( n220 , n25 , n37 );
not ( n221 , n220 );
not ( n222 , n221 );
not ( n223 , n222 );
not ( n224 , n185 );
not ( n225 , n224 );
or ( n226 , n223 , n225 );
not ( n227 , n135 );
not ( n228 , n227 );
nand ( n229 , n226 , n228 );
or ( n230 , n33 , n229 );
not ( n231 , n32 );
not ( n232 , n37 );
or ( n233 , n232 , n26 );
not ( n234 , n25 );
nand ( n235 , n233 , n234 );
and ( n236 , n231 , n235 );
not ( n237 , n236 );
not ( n238 , n193 );
nand ( n239 , n238 , n187 , n168 , n182 );
not ( n240 , n239 );
or ( n241 , n237 , n240 );
nor ( n242 , n185 , n32 );
nor ( n243 , n25 , n37 );
nand ( n244 , n136 , n242 , n243 );
not ( n245 , n244 );
not ( n246 , n32 );
and ( n247 , n246 , n227 );
nor ( n248 , n245 , n247 );
nand ( n249 , n241 , n248 );
nand ( n250 , n230 , n249 );
nand ( n251 , n212 , n219 , n250 );
not ( n252 , n251 );
or ( n253 , n155 , n252 );
not ( n254 , n35 );
nor ( n255 , n254 , n32 );
not ( n256 , n255 );
and ( n257 , n256 , n211 );
not ( n258 , n122 );
not ( n259 , n258 );
nand ( n260 , n26 , n259 );
not ( n261 , n26 );
not ( n262 , n185 );
not ( n263 , n262 );
nand ( n264 , n261 , n263 );
nand ( n265 , n260 , n234 , n264 );
not ( n266 , n265 );
and ( n267 , n266 , n256 );
nor ( n268 , n257 , n267 );
nand ( n269 , n253 , n268 );
not ( n270 , n269 );
not ( n271 , n270 );
or ( n272 , n154 , n271 );
not ( n273 , n23 );
and ( n274 , n22 , n273 );
not ( n275 , n274 );
buf ( n276 , n275 );
not ( n277 , n276 );
not ( n278 , n277 );
not ( n279 , n278 );
not ( n280 , n279 );
buf ( n281 , n280 );
nand ( n282 , n272 , n281 );
nand ( n283 , n147 , n282 );
nand ( n284 , n140 , n283 );
nand ( n285 , n82 , n99 , n18 , n284 );
buf ( n286 , n90 );
not ( n287 , n286 );
not ( n288 , n287 );
not ( n289 , n288 );
not ( n290 , n289 );
not ( n291 , n290 );
not ( n292 , n291 );
not ( n293 , n18 );
or ( n294 , n293 , n19 );
not ( n295 , n96 );
nor ( n296 , n294 , n295 );
not ( n297 , n24 );
nor ( n298 , n297 , n31 );
or ( n299 , n100 , n298 );
and ( n300 , n299 , n105 , n138 );
nand ( n301 , n300 , n283 );
nand ( n302 , n292 , n296 , n82 , n301 );
not ( n303 , n19 );
not ( n304 , n14 );
nand ( n305 , n16 , n304 );
and ( n306 , n303 , n305 );
not ( n307 , n18 );
or ( n308 , n307 , n20 );
not ( n309 , n308 );
not ( n310 , n23 );
nor ( n311 , n310 , n298 );
not ( n312 , n311 );
nand ( n313 , n23 , n312 );
nand ( n314 , n22 , n313 );
and ( n315 , n87 , n314 );
not ( n316 , n22 );
and ( n317 , n316 , n86 );
nor ( n318 , n315 , n317 , n17 );
not ( n319 , n318 );
not ( n320 , n23 );
not ( n321 , n22 );
nor ( n322 , n28 , n31 );
not ( n323 , n322 );
nand ( n324 , n321 , n323 );
nand ( n325 , n320 , n324 );
nand ( n326 , n299 , n325 );
and ( n327 , n326 , n87 );
nand ( n328 , n100 , n325 );
and ( n329 , n86 , n328 );
nor ( n330 , n327 , n329 );
nor ( n331 , n15 , n330 );
nand ( n332 , n17 , n331 );
and ( n333 , n319 , n332 );
not ( n334 , n333 );
nand ( n335 , n306 , n80 , n309 , n334 );
buf ( n336 , n146 );
not ( n337 , n336 );
and ( n338 , n234 , n224 );
nor ( n339 , n25 , n109 );
not ( n340 , n339 );
nor ( n341 , n338 , n26 , n340 );
not ( n342 , n341 );
not ( n343 , n342 );
buf ( n344 , n249 );
not ( n345 , n344 );
and ( n346 , n343 , n345 );
nor ( n347 , n346 , n279 );
or ( n348 , n25 , n26 );
not ( n349 , n348 );
not ( n350 , n349 );
not ( n351 , n350 );
nand ( n352 , n32 , n351 , n224 );
nand ( n353 , n234 , n258 );
and ( n354 , n353 , n26 , n339 );
nor ( n355 , n32 , n23 , n31 );
nor ( n356 , n354 , n355 );
or ( n357 , n356 , n344 );
nand ( n358 , n248 , n149 , n228 );
buf ( n359 , n195 );
or ( n360 , n358 , n359 );
nand ( n361 , n360 , n276 );
not ( n362 , n361 );
nand ( n363 , n357 , n362 );
nand ( n364 , n352 , n363 );
and ( n365 , n347 , n364 );
not ( n366 , n365 );
and ( n367 , n337 , n366 );
nor ( n368 , n367 , n139 );
and ( n369 , n14 , n368 );
not ( n370 , n14 );
nor ( n371 , n232 , n25 );
nand ( n372 , n242 , n371 , n136 );
not ( n373 , n247 );
nand ( n374 , n372 , n373 );
not ( n375 , n374 );
buf ( n376 , n375 );
buf ( n377 , n376 );
not ( n378 , n32 );
nor ( n379 , n26 , n37 );
not ( n380 , n379 );
nand ( n381 , n234 , n380 );
and ( n382 , n378 , n381 );
not ( n383 , n187 );
nor ( n384 , n34 , n36 );
not ( n385 , n384 );
nand ( n386 , n385 , n175 );
not ( n387 , n386 );
not ( n388 , n387 );
not ( n389 , n166 );
buf ( n390 , n389 );
not ( n391 , n30 );
nand ( n392 , n36 , n391 );
not ( n393 , n392 );
nand ( n394 , n388 , n390 , n393 );
not ( n395 , n394 );
nor ( n396 , n383 , n395 );
not ( n397 , n387 );
nand ( n398 , n181 , n397 );
not ( n399 , n167 );
and ( n400 , n398 , n399 );
nand ( n401 , n396 , n400 );
buf ( n402 , n401 );
nand ( n403 , n382 , n402 );
nand ( n404 , n377 , n341 , n403 );
not ( n405 , n148 );
nand ( n406 , n405 , n228 );
nor ( n407 , n374 , n406 );
buf ( n408 , n407 );
not ( n409 , n402 );
and ( n410 , n408 , n409 );
not ( n411 , n276 );
nor ( n412 , n410 , n411 );
not ( n413 , n356 );
nand ( n414 , n413 , n376 , n403 );
nand ( n415 , n412 , n414 );
and ( n416 , n352 , n415 );
not ( n417 , n280 );
nor ( n418 , n416 , n417 );
nand ( n419 , n404 , n418 );
and ( n420 , n337 , n419 );
nor ( n421 , n420 , n139 );
and ( n422 , n370 , n421 );
not ( n423 , n19 );
not ( n424 , n16 );
nand ( n425 , n15 , n17 );
not ( n426 , n425 );
nand ( n427 , n423 , n424 , n426 );
not ( n428 , n427 );
not ( n429 , n428 );
not ( n430 , n429 );
buf ( n431 , n430 );
not ( n432 , n431 );
not ( n433 , n432 );
not ( n434 , n433 );
not ( n435 , n434 );
not ( n436 , n435 );
not ( n437 , n436 );
not ( n438 , n437 );
nor ( n439 , n369 , n422 , n438 );
nor ( n440 , n20 , n90 );
not ( n441 , n18 );
nor ( n442 , n441 , n81 );
nand ( n443 , n439 , n440 , n442 );
and ( n444 , n285 , n302 , n335 , n443 );
not ( n445 , n41 );
not ( n446 , n14 );
not ( n447 , n426 );
buf ( n448 , n447 );
not ( n449 , n448 );
and ( n450 , n446 , n449 );
not ( n451 , n19 );
not ( n452 , n20 );
and ( n453 , n451 , n452 );
and ( n454 , n16 , n453 );
nand ( n455 , n450 , n454 );
nor ( n456 , n40 , n455 );
nand ( n457 , n445 , n456 );
not ( n458 , n457 );
not ( n459 , n147 );
not ( n460 , n459 );
not ( n461 , n153 );
not ( n462 , n461 );
not ( n463 , n462 );
not ( n464 , n217 );
nand ( n465 , n232 , n214 );
nor ( n466 , n33 , n465 );
and ( n467 , n464 , n466 );
not ( n468 , n467 );
not ( n469 , n382 );
not ( n470 , n401 );
or ( n471 , n469 , n470 );
nand ( n472 , n471 , n375 );
not ( n473 , n33 );
not ( n474 , n37 );
nor ( n475 , n474 , n25 );
not ( n476 , n475 );
not ( n477 , n476 );
not ( n478 , n477 );
not ( n479 , n181 );
or ( n480 , n478 , n479 );
nand ( n481 , n480 , n228 );
not ( n482 , n481 );
nand ( n483 , n473 , n482 );
nand ( n484 , n472 , n483 );
nand ( n485 , n468 , n484 );
not ( n486 , n32 );
not ( n487 , n161 );
not ( n488 , n487 );
not ( n489 , n401 );
or ( n490 , n488 , n489 );
nand ( n491 , n490 , n210 );
nand ( n492 , n486 , n491 );
not ( n493 , n492 );
nor ( n494 , n485 , n493 );
not ( n495 , n35 );
nor ( n496 , n494 , n495 );
not ( n497 , n256 );
not ( n498 , n491 );
or ( n499 , n497 , n498 );
not ( n500 , n267 );
nand ( n501 , n499 , n500 );
nor ( n502 , n496 , n501 );
not ( n503 , n502 );
or ( n504 , n463 , n503 );
buf ( n505 , n281 );
nand ( n506 , n504 , n505 );
nand ( n507 , n460 , n506 );
nand ( n508 , n300 , n507 );
and ( n509 , n442 , n458 , n508 );
nand ( n510 , n140 , n507 );
nor ( n511 , n90 , n455 );
and ( n512 , n510 , n442 , n511 );
nor ( n513 , n509 , n512 );
not ( n514 , n20 );
and ( n515 , n19 , n514 );
not ( n516 , n515 );
not ( n517 , n17 );
nor ( n518 , n517 , n16 );
not ( n519 , n14 );
and ( n520 , n518 , n15 , n519 );
not ( n521 , n520 );
nor ( n522 , n516 , n521 );
not ( n523 , n522 );
not ( n524 , n147 );
not ( n525 , n524 );
not ( n526 , n525 );
nor ( n527 , n523 , n526 );
not ( n528 , n462 );
not ( n529 , n35 );
not ( n530 , n33 );
nor ( n531 , n465 , n530 );
and ( n532 , n531 , n218 );
not ( n533 , n532 );
not ( n534 , n202 );
not ( n535 , n534 );
not ( n536 , n401 );
or ( n537 , n535 , n536 );
not ( n538 , n161 );
nand ( n539 , n209 , n538 );
buf ( n540 , n539 );
nand ( n541 , n537 , n540 );
not ( n542 , n32 );
nand ( n543 , n541 , n542 );
not ( n544 , n33 );
or ( n545 , n481 , n544 );
nand ( n546 , n545 , n472 );
nand ( n547 , n533 , n543 , n546 );
nand ( n548 , n529 , n547 );
or ( n549 , n32 , n35 );
not ( n550 , n549 );
not ( n551 , n550 );
not ( n552 , n551 );
buf ( n553 , n552 );
not ( n554 , n553 );
and ( n555 , n554 , n541 );
or ( n556 , n265 , n552 );
not ( n557 , n556 );
nor ( n558 , n555 , n557 );
nand ( n559 , n548 , n558 );
not ( n560 , n559 );
not ( n561 , n560 );
or ( n562 , n528 , n561 );
buf ( n563 , n281 );
nand ( n564 , n562 , n563 );
not ( n565 , n564 );
not ( n566 , n565 );
and ( n567 , n527 , n566 );
buf ( n568 , n95 );
buf ( n569 , n568 );
and ( n570 , n515 , n569 );
not ( n571 , n570 );
not ( n572 , n524 );
not ( n573 , n572 );
nor ( n574 , n571 , n573 );
nand ( n575 , n25 , n218 );
nor ( n576 , n150 , n266 );
and ( n577 , n575 , n576 );
nor ( n578 , n577 , n411 );
not ( n579 , n578 );
and ( n580 , n574 , n579 );
nor ( n581 , n567 , n580 );
not ( n582 , n20 );
and ( n583 , n19 , n520 );
and ( n584 , n582 , n583 );
not ( n585 , n584 );
nor ( n586 , n585 , n300 );
not ( n587 , n586 );
and ( n588 , n14 , n15 );
not ( n589 , n16 );
and ( n590 , n588 , n589 , n17 );
nand ( n591 , n515 , n590 );
nor ( n592 , n591 , n526 );
not ( n593 , n153 );
not ( n594 , n33 );
or ( n595 , n229 , n594 );
nand ( n596 , n249 , n595 );
not ( n597 , n534 );
not ( n598 , n239 );
or ( n599 , n597 , n598 );
nand ( n600 , n599 , n539 );
not ( n601 , n32 );
nand ( n602 , n600 , n601 );
not ( n603 , n26 );
not ( n604 , n32 );
nand ( n605 , n604 , n37 );
not ( n606 , n605 );
nand ( n607 , n33 , n603 , n606 );
or ( n608 , n217 , n607 );
nand ( n609 , n596 , n602 , n608 );
not ( n610 , n35 );
nand ( n611 , n609 , n610 );
not ( n612 , n556 );
not ( n613 , n612 );
not ( n614 , n553 );
nand ( n615 , n600 , n614 );
buf ( n616 , n615 );
nand ( n617 , n611 , n613 , n616 );
not ( n618 , n617 );
not ( n619 , n618 );
or ( n620 , n593 , n619 );
nand ( n621 , n620 , n505 );
and ( n622 , n592 , n621 );
not ( n623 , n515 );
not ( n624 , n623 );
not ( n625 , n624 );
not ( n626 , n625 );
not ( n627 , n626 );
buf ( n628 , n627 );
not ( n629 , n628 );
not ( n630 , n629 );
not ( n631 , n569 );
not ( n632 , n590 );
and ( n633 , n631 , n632 );
nor ( n634 , n630 , n633 , n300 );
nor ( n635 , n622 , n634 );
nand ( n636 , n581 , n587 , n635 );
not ( n637 , n292 );
not ( n638 , n637 );
nand ( n639 , n636 , n638 , n442 );
not ( n640 , n19 );
nand ( n641 , n640 , n20 );
not ( n642 , n641 );
not ( n643 , n642 );
not ( n644 , n643 );
not ( n645 , n644 );
not ( n646 , n645 );
nand ( n647 , n646 , n96 );
nor ( n648 , n40 , n647 );
not ( n649 , n153 );
not ( n650 , n35 );
not ( n651 , n487 );
and ( n652 , n164 , n34 );
buf ( n653 , n652 );
nor ( n654 , n653 , n193 );
not ( n655 , n179 );
and ( n656 , n655 , n262 );
nor ( n657 , n656 , n167 );
nand ( n658 , n654 , n657 );
not ( n659 , n658 );
or ( n660 , n651 , n659 );
nand ( n661 , n201 , n206 );
not ( n662 , n661 );
not ( n663 , n662 );
nand ( n664 , n660 , n663 );
not ( n665 , n32 );
and ( n666 , n664 , n665 );
not ( n667 , n206 );
nor ( n668 , n667 , n215 );
nor ( n669 , n666 , n668 );
not ( n670 , n236 );
not ( n671 , n658 );
or ( n672 , n670 , n671 );
nand ( n673 , n672 , n248 );
nand ( n674 , n230 , n673 );
nand ( n675 , n669 , n674 );
not ( n676 , n675 );
or ( n677 , n650 , n676 );
not ( n678 , n664 );
not ( n679 , n678 );
and ( n680 , n256 , n679 );
nor ( n681 , n680 , n267 );
nand ( n682 , n677 , n681 );
not ( n683 , n682 );
not ( n684 , n683 );
or ( n685 , n649 , n684 );
nand ( n686 , n685 , n281 );
nand ( n687 , n147 , n686 );
nand ( n688 , n140 , n687 );
and ( n689 , n648 , n688 );
not ( n690 , n20 );
not ( n691 , n15 );
nand ( n692 , n691 , n17 );
not ( n693 , n692 );
nand ( n694 , n40 , n693 , n326 );
not ( n695 , n40 );
not ( n696 , n17 );
not ( n697 , n23 );
not ( n698 , n697 );
not ( n699 , n322 );
or ( n700 , n698 , n699 );
not ( n701 , n22 );
nand ( n702 , n700 , n701 );
and ( n703 , n92 , n702 );
not ( n704 , n703 );
nor ( n705 , n696 , n704 );
and ( n706 , n695 , n705 );
and ( n707 , n40 , n314 );
not ( n708 , n22 );
not ( n709 , n40 );
and ( n710 , n708 , n709 );
nor ( n711 , n707 , n710 , n17 );
nor ( n712 , n706 , n711 );
and ( n713 , n694 , n712 );
nor ( n714 , n690 , n713 );
nor ( n715 , n689 , n714 );
not ( n716 , n647 );
nand ( n717 , n40 , n716 );
not ( n718 , n717 );
nand ( n719 , n300 , n687 );
not ( n720 , n719 );
not ( n721 , n720 );
and ( n722 , n718 , n721 );
not ( n723 , n14 );
and ( n724 , n723 , n95 );
nand ( n725 , n644 , n724 );
nor ( n726 , n40 , n725 );
not ( n727 , n726 );
not ( n728 , n35 );
not ( n729 , n483 );
not ( n730 , n374 );
not ( n731 , n652 );
nand ( n732 , n398 , n394 , n168 , n731 );
nand ( n733 , n732 , n382 );
nand ( n734 , n730 , n733 );
not ( n735 , n734 );
or ( n736 , n729 , n735 );
not ( n737 , n667 );
not ( n738 , n466 );
not ( n739 , n738 );
and ( n740 , n737 , n739 );
not ( n741 , n487 );
not ( n742 , n732 );
or ( n743 , n741 , n742 );
not ( n744 , n662 );
nand ( n745 , n743 , n744 );
not ( n746 , n32 );
and ( n747 , n745 , n746 );
nor ( n748 , n740 , n747 );
nand ( n749 , n736 , n748 );
not ( n750 , n749 );
or ( n751 , n728 , n750 );
and ( n752 , n256 , n745 );
nor ( n753 , n752 , n267 );
nand ( n754 , n751 , n753 );
or ( n755 , n461 , n754 );
nand ( n756 , n755 , n281 );
nand ( n757 , n337 , n756 );
nand ( n758 , n140 , n757 );
not ( n759 , n758 );
nor ( n760 , n727 , n759 );
nor ( n761 , n722 , n760 );
not ( n762 , n40 );
not ( n763 , n20 );
and ( n764 , n19 , n590 );
nand ( n765 , n763 , n764 );
not ( n766 , n765 );
not ( n767 , n766 );
not ( n768 , n336 );
not ( n769 , n768 );
not ( n770 , n621 );
or ( n771 , n769 , n770 );
nand ( n772 , n771 , n140 );
not ( n773 , n772 );
or ( n774 , n767 , n773 );
not ( n775 , n572 );
not ( n776 , n564 );
or ( n777 , n775 , n776 );
nand ( n778 , n777 , n140 );
and ( n779 , n584 , n778 );
not ( n780 , n20 );
and ( n781 , n19 , n569 );
and ( n782 , n780 , n781 );
or ( n783 , n146 , n578 );
nand ( n784 , n783 , n140 );
and ( n785 , n782 , n784 );
nor ( n786 , n779 , n785 );
nand ( n787 , n774 , n786 );
and ( n788 , n762 , n787 );
nand ( n789 , n453 , n724 );
nor ( n790 , n40 , n789 );
and ( n791 , n790 , n510 );
nor ( n792 , n788 , n791 );
and ( n793 , n40 , n636 );
nand ( n794 , n20 , n40 );
or ( n795 , n14 , n427 );
nor ( n796 , n795 , n143 );
nand ( n797 , n377 , n341 , n733 );
buf ( n798 , n732 );
not ( n799 , n798 );
and ( n800 , n799 , n407 );
not ( n801 , n276 );
nor ( n802 , n800 , n801 );
not ( n803 , n356 );
nand ( n804 , n803 , n375 , n733 );
nand ( n805 , n802 , n804 );
nand ( n806 , n352 , n805 );
and ( n807 , n797 , n280 , n806 );
not ( n808 , n807 );
nand ( n809 , n796 , n808 );
not ( n810 , n809 );
not ( n811 , n300 );
nand ( n812 , n433 , n811 );
not ( n813 , n812 );
not ( n814 , n673 );
and ( n815 , n341 , n814 );
nor ( n816 , n815 , n279 );
not ( n817 , n356 );
nand ( n818 , n817 , n814 );
not ( n819 , n358 );
not ( n820 , n653 );
and ( n821 , n238 , n820 , n168 , n182 );
not ( n822 , n821 );
not ( n823 , n822 );
nand ( n824 , n819 , n823 );
nand ( n825 , n818 , n278 , n824 );
nand ( n826 , n352 , n825 );
and ( n827 , n816 , n826 );
not ( n828 , n428 );
not ( n829 , n14 );
nor ( n830 , n828 , n829 );
nand ( n831 , n830 , n144 );
nor ( n832 , n827 , n831 );
nor ( n833 , n810 , n813 , n832 );
nor ( n834 , n794 , n833 );
nor ( n835 , n793 , n834 );
nand ( n836 , n715 , n761 , n792 , n835 );
not ( n837 , n40 );
nor ( n838 , n837 , n789 );
and ( n839 , n838 , n508 );
not ( n840 , n40 );
not ( n841 , n453 );
nor ( n842 , n841 , n295 );
not ( n843 , n842 );
nor ( n844 , n840 , n843 );
not ( n845 , n844 );
not ( n846 , n301 );
or ( n847 , n845 , n846 );
nor ( n848 , n40 , n843 );
nand ( n849 , n848 , n284 );
nand ( n850 , n847 , n849 );
nor ( n851 , n20 , n713 );
nor ( n852 , n839 , n850 , n851 );
nor ( n853 , n20 , n40 );
and ( n854 , n853 , n439 );
not ( n855 , n40 );
nor ( n856 , n855 , n20 );
not ( n857 , n419 );
buf ( n858 , n857 );
not ( n859 , n858 );
and ( n860 , n796 , n859 );
or ( n861 , n831 , n365 );
nand ( n862 , n861 , n812 );
nor ( n863 , n860 , n862 );
not ( n864 , n863 );
and ( n865 , n856 , n864 );
nor ( n866 , n854 , n865 );
not ( n867 , n40 );
nand ( n868 , n20 , n867 );
not ( n869 , n868 );
nand ( n870 , n431 , n139 );
not ( n871 , n832 );
nand ( n872 , n809 , n870 , n871 );
and ( n873 , n869 , n872 );
not ( n874 , n40 );
nor ( n875 , n874 , n725 );
and ( n876 , n300 , n757 );
not ( n877 , n876 );
and ( n878 , n875 , n877 );
nor ( n879 , n873 , n878 );
not ( n880 , n40 );
not ( n881 , n462 );
not ( n882 , n534 );
not ( n883 , n732 );
or ( n884 , n882 , n883 );
not ( n885 , n206 );
or ( n886 , n159 , n885 );
nand ( n887 , n884 , n886 );
not ( n888 , n887 );
nor ( n889 , n888 , n553 );
not ( n890 , n889 );
not ( n891 , n35 );
not ( n892 , n32 );
nand ( n893 , n887 , n892 );
nand ( n894 , n734 , n545 );
not ( n895 , n531 );
or ( n896 , n895 , n667 );
nand ( n897 , n893 , n894 , n896 );
nand ( n898 , n891 , n897 );
not ( n899 , n612 );
nand ( n900 , n890 , n898 , n899 );
not ( n901 , n900 );
not ( n902 , n901 );
or ( n903 , n881 , n902 );
nand ( n904 , n903 , n563 );
nand ( n905 , n337 , n904 );
nand ( n906 , n140 , n905 );
not ( n907 , n906 );
and ( n908 , n19 , n20 );
and ( n909 , n908 , n520 );
not ( n910 , n909 );
or ( n911 , n907 , n910 );
not ( n912 , n908 );
or ( n913 , n912 , n632 );
not ( n914 , n913 );
not ( n915 , n461 );
not ( n916 , n915 );
not ( n917 , n35 );
nand ( n918 , n673 , n595 );
not ( n919 , n32 );
not ( n920 , n202 );
not ( n921 , n920 );
not ( n922 , n658 );
or ( n923 , n921 , n922 );
nand ( n924 , n923 , n886 );
nand ( n925 , n919 , n924 );
not ( n926 , n667 );
not ( n927 , n607 );
nand ( n928 , n926 , n927 );
nand ( n929 , n918 , n925 , n928 );
nand ( n930 , n917 , n929 );
nand ( n931 , n614 , n924 );
nand ( n932 , n930 , n931 , n613 );
not ( n933 , n932 );
not ( n934 , n933 );
or ( n935 , n916 , n934 );
nand ( n936 , n935 , n505 );
not ( n937 , n936 );
not ( n938 , n768 );
or ( n939 , n937 , n938 );
nand ( n940 , n939 , n140 );
and ( n941 , n914 , n940 );
and ( n942 , n908 , n568 );
not ( n943 , n145 );
not ( n944 , n926 );
nor ( n945 , n234 , n944 );
not ( n946 , n945 );
nand ( n947 , n946 , n576 );
and ( n948 , n280 , n947 );
or ( n949 , n943 , n948 );
nand ( n950 , n949 , n140 );
and ( n951 , n942 , n950 );
nor ( n952 , n941 , n951 );
nand ( n953 , n911 , n952 );
and ( n954 , n880 , n953 );
nand ( n955 , n909 , n525 );
not ( n956 , n904 );
not ( n957 , n956 );
not ( n958 , n957 );
or ( n959 , n955 , n958 );
not ( n960 , n936 );
nand ( n961 , n914 , n147 );
or ( n962 , n960 , n961 );
not ( n963 , n942 );
not ( n964 , n145 );
nor ( n965 , n963 , n964 );
not ( n966 , n948 );
and ( n967 , n965 , n966 );
and ( n968 , n914 , n811 );
nor ( n969 , n967 , n968 );
buf ( n970 , n631 );
buf ( n971 , n970 );
buf ( n972 , n971 );
not ( n973 , n972 );
or ( n974 , n973 , n520 );
nor ( n975 , n912 , n300 );
nand ( n976 , n974 , n975 );
nand ( n977 , n962 , n969 , n976 );
not ( n978 , n977 );
nand ( n979 , n959 , n978 );
and ( n980 , n40 , n979 );
nor ( n981 , n954 , n980 );
nand ( n982 , n852 , n866 , n879 , n981 );
or ( n983 , n836 , n982 );
not ( n984 , n18 );
nor ( n985 , n12 , n78 );
nand ( n986 , n13 , n985 );
not ( n987 , n986 );
not ( n988 , n987 );
nor ( n989 , n984 , n988 );
nand ( n990 , n983 , n989 );
nand ( n991 , n444 , n513 , n639 , n990 );
not ( n992 , n2 );
and ( n993 , n12 , n992 );
and ( n994 , n11 , n993 );
not ( n995 , n994 );
not ( n996 , n995 );
not ( n997 , n35 );
not ( n998 , n31 );
not ( n999 , n23 );
nand ( n1000 , n26 , n32 );
and ( n1001 , n998 , n999 , n1000 );
nand ( n1002 , n997 , n32 , n1001 );
not ( n1003 , n1002 );
not ( n1004 , n26 );
not ( n1005 , n32 );
nor ( n1006 , n1005 , n33 );
and ( n1007 , n1004 , n1006 );
buf ( n1008 , n1007 );
nand ( n1009 , n209 , n1008 );
not ( n1010 , n32 );
nor ( n1011 , n135 , n1010 );
not ( n1012 , n1011 );
and ( n1013 , n1009 , n1012 );
not ( n1014 , n1013 );
not ( n1015 , n1014 );
not ( n1016 , n359 );
buf ( n1017 , n1016 );
buf ( n1018 , n1017 );
and ( n1019 , n1003 , n1015 , n1018 );
buf ( n1020 , n211 );
nand ( n1021 , n32 , n110 );
nor ( n1022 , n35 , n1021 );
and ( n1023 , n1022 , n1009 );
not ( n1024 , n26 );
and ( n1025 , n33 , n1024 );
nand ( n1026 , n32 , n1025 );
not ( n1027 , n1012 );
not ( n1028 , n1027 );
nand ( n1029 , n1023 , n1026 , n1028 );
not ( n1030 , n359 );
nand ( n1031 , n1023 , n1028 , n1030 );
and ( n1032 , n1029 , n1031 );
or ( n1033 , n1020 , n1032 );
nor ( n1034 , n1025 , n1002 );
and ( n1035 , n1034 , n1013 );
nor ( n1036 , n1035 , n411 );
nand ( n1037 , n1033 , n1036 );
nor ( n1038 , n1019 , n1037 );
not ( n1039 , n1020 );
not ( n1040 , n1039 );
not ( n1041 , n1015 );
buf ( n1042 , n1030 );
not ( n1043 , n1042 );
nor ( n1044 , n1040 , n1041 , n1043 );
not ( n1045 , n35 );
not ( n1046 , n23 );
and ( n1047 , n1045 , n1046 , n998 );
nand ( n1048 , n1044 , n1047 , n270 );
nand ( n1049 , n1038 , n1048 );
not ( n1050 , n23 );
and ( n1051 , n32 , n1050 );
and ( n1052 , n998 , n1051 );
nor ( n1053 , n26 , n33 );
not ( n1054 , n1053 );
nand ( n1055 , n32 , n1054 );
nand ( n1056 , n1015 , n1052 , n1055 );
not ( n1057 , n1056 );
not ( n1058 , n1020 );
nand ( n1059 , n1052 , n1058 , n1015 , n1017 );
not ( n1060 , n1059 );
or ( n1061 , n1057 , n1060 );
not ( n1062 , n251 );
nand ( n1063 , n1061 , n1062 );
and ( n1064 , n1001 , n1009 );
buf ( n1065 , n1027 );
not ( n1066 , n1065 );
not ( n1067 , n1066 );
not ( n1068 , n1067 );
and ( n1069 , n1064 , n1026 , n1068 );
nand ( n1070 , n270 , n1062 , n1069 );
nand ( n1071 , n1063 , n1070 );
nor ( n1072 , n1049 , n1071 );
not ( n1073 , n1020 );
not ( n1074 , n23 );
nand ( n1075 , n32 , n33 );
not ( n1076 , n1075 );
not ( n1077 , n26 );
and ( n1078 , n1076 , n1077 );
not ( n1079 , n1078 );
nand ( n1080 , n1074 , n1079 , n1009 );
not ( n1081 , n1080 );
nand ( n1082 , n1081 , n998 , n1028 );
not ( n1083 , n1082 );
and ( n1084 , n1073 , n1083 , n1062 );
not ( n1085 , n1055 );
not ( n1086 , n1047 );
nor ( n1087 , n1014 , n1085 , n1086 );
nor ( n1088 , n1084 , n1087 );
or ( n1089 , n269 , n1088 );
not ( n1090 , n1040 );
not ( n1091 , n32 );
nor ( n1092 , n1082 , n1091 );
nand ( n1093 , n1090 , n1092 , n1062 );
nor ( n1094 , n26 , n109 );
and ( n1095 , n32 , n1094 );
and ( n1096 , n1095 , n1009 );
and ( n1097 , n1096 , n1017 );
not ( n1098 , n1065 );
and ( n1099 , n1098 , n212 );
nand ( n1100 , n1097 , n219 , n1099 , n250 );
nand ( n1101 , n1089 , n1093 , n1100 );
not ( n1102 , n1068 );
not ( n1103 , n1102 );
not ( n1104 , n1000 );
not ( n1105 , n1104 );
nand ( n1106 , n1009 , n1105 , n1047 );
nor ( n1107 , n1106 , n1043 );
nand ( n1108 , n270 , n1103 , n1107 );
not ( n1109 , n35 );
nand ( n1110 , n1109 , n1083 );
not ( n1111 , n1110 );
nand ( n1112 , n1111 , n1073 );
not ( n1113 , n1112 );
not ( n1114 , n219 );
not ( n1115 , n359 );
buf ( n1116 , n1115 );
not ( n1117 , n1116 );
nor ( n1118 , n1114 , n1117 );
nand ( n1119 , n1118 , n1064 , n1099 , n250 );
not ( n1120 , n1119 );
or ( n1121 , n1113 , n1120 );
nand ( n1122 , n1121 , n270 );
and ( n1123 , n1039 , n1015 , n268 );
nor ( n1124 , n150 , n359 );
nand ( n1125 , n1123 , n1124 , n1062 );
nand ( n1126 , n1108 , n1122 , n1125 );
nor ( n1127 , n1101 , n1126 );
nand ( n1128 , n1072 , n1127 );
not ( n1129 , n525 );
not ( n1130 , n1129 );
nand ( n1131 , n1128 , n1130 );
nand ( n1132 , n1131 , n140 );
not ( n1133 , n20 );
nor ( n1134 , n18 , n19 );
not ( n1135 , n1134 );
nor ( n1136 , n1135 , n295 );
and ( n1137 , n1133 , n1136 );
and ( n1138 , n1132 , n1137 );
not ( n1139 , n20 );
not ( n1140 , n18 );
nand ( n1141 , n1140 , n430 );
nor ( n1142 , n14 , n1141 );
nand ( n1143 , n1139 , n1142 );
not ( n1144 , n1143 );
not ( n1145 , n415 );
or ( n1146 , n459 , n1145 );
nand ( n1147 , n1146 , n140 );
and ( n1148 , n1144 , n1147 );
nor ( n1149 , n1138 , n1148 );
not ( n1150 , n502 );
not ( n1151 , n162 );
not ( n1152 , n1151 );
not ( n1153 , n1152 );
not ( n1154 , n402 );
or ( n1155 , n1153 , n1154 );
nand ( n1156 , n1155 , n210 );
or ( n1157 , n1110 , n1156 );
not ( n1158 , n409 );
not ( n1159 , n1158 );
not ( n1160 , n1065 );
and ( n1161 , n1160 , n492 );
not ( n1162 , n485 );
nand ( n1163 , n1064 , n1159 , n1161 , n1162 );
nand ( n1164 , n1157 , n1163 );
not ( n1165 , n1164 );
or ( n1166 , n1150 , n1165 );
nor ( n1167 , n1102 , n1106 , n501 );
not ( n1168 , n496 );
not ( n1169 , n1159 );
not ( n1170 , n1169 );
and ( n1171 , n1167 , n1168 , n1170 );
buf ( n1172 , n491 );
nor ( n1173 , n501 , n152 , n1172 );
not ( n1174 , n1014 );
and ( n1175 , n1174 , n409 );
and ( n1176 , n1173 , n1175 , n494 );
nor ( n1177 , n1171 , n1176 );
nand ( n1178 , n1166 , n1177 );
not ( n1179 , n502 );
not ( n1180 , n1087 );
not ( n1181 , n467 );
not ( n1182 , n484 );
nor ( n1183 , n493 , n1156 , n1182 );
nand ( n1184 , n1181 , n1183 , n1083 );
nand ( n1185 , n1180 , n1184 );
not ( n1186 , n1185 );
or ( n1187 , n1179 , n1186 );
not ( n1188 , n1161 );
nor ( n1189 , n1188 , n467 , n1182 );
and ( n1190 , n1096 , n1189 , n1170 );
not ( n1191 , n1156 );
not ( n1192 , n1182 );
nand ( n1193 , n1191 , n1092 , n1192 );
nor ( n1194 , n1193 , n467 , n493 );
nor ( n1195 , n1190 , n1194 );
nand ( n1196 , n1187 , n1195 );
nor ( n1197 , n1178 , n1196 );
buf ( n1198 , n1172 );
nor ( n1199 , n1086 , n1198 );
and ( n1200 , n1199 , n1175 , n502 );
and ( n1201 , n1068 , n1023 , n1159 );
not ( n1202 , n1029 );
nor ( n1203 , n1201 , n1202 );
or ( n1204 , n1203 , n1198 );
nand ( n1205 , n1003 , n1175 );
nand ( n1206 , n1204 , n1205 , n1036 );
nor ( n1207 , n1200 , n1206 );
not ( n1208 , n494 );
not ( n1209 , n1208 );
and ( n1210 , n1069 , n1209 , n502 );
not ( n1211 , n1198 );
and ( n1212 , n1211 , n1052 , n1175 );
not ( n1213 , n1056 );
nor ( n1214 , n1212 , n1213 );
nor ( n1215 , n1214 , n1208 );
nor ( n1216 , n1210 , n1215 );
nand ( n1217 , n1197 , n1207 , n1216 );
not ( n1218 , n1217 );
not ( n1219 , n1218 );
nand ( n1220 , n1219 , n1130 );
nand ( n1221 , n140 , n1220 );
nand ( n1222 , n1134 , n724 );
nor ( n1223 , n20 , n1222 );
nand ( n1224 , n1221 , n1223 );
not ( n1225 , n768 );
not ( n1226 , n1225 );
not ( n1227 , n1011 );
nand ( n1228 , n206 , n1007 );
and ( n1229 , n1227 , n1228 );
buf ( n1230 , n1229 );
and ( n1231 , n1034 , n1230 );
nor ( n1232 , n1231 , n279 );
buf ( n1233 , n1230 );
not ( n1234 , n1233 );
not ( n1235 , n1234 );
not ( n1236 , n798 );
buf ( n1237 , n1236 );
nand ( n1238 , n1235 , n1003 , n1237 );
buf ( n1239 , n1079 );
not ( n1240 , n1239 );
nand ( n1241 , n1022 , n1229 );
nor ( n1242 , n1240 , n1241 );
not ( n1243 , n745 );
and ( n1244 , n1242 , n1243 );
not ( n1245 , n1241 );
not ( n1246 , n798 );
and ( n1247 , n744 , n1246 );
and ( n1248 , n1245 , n1247 );
nor ( n1249 , n1244 , n1248 );
and ( n1250 , n1232 , n1238 , n1249 );
not ( n1251 , n1052 );
buf ( n1252 , n1229 );
and ( n1253 , n1055 , n1252 );
not ( n1254 , n1253 );
nor ( n1255 , n1251 , n1254 );
not ( n1256 , n1255 );
not ( n1257 , n749 );
not ( n1258 , n1257 );
or ( n1259 , n1256 , n1258 );
buf ( n1260 , n1230 );
not ( n1261 , n1095 );
nor ( n1262 , n1261 , n798 );
nand ( n1263 , n1260 , n1262 , n1257 );
nand ( n1264 , n1259 , n1263 );
not ( n1265 , n32 );
not ( n1266 , n23 );
nand ( n1267 , n1266 , n1252 );
nor ( n1268 , n1265 , n31 , n1267 );
nand ( n1269 , n1257 , n1247 , n1268 );
and ( n1270 , n1230 , n1239 , n1052 );
nand ( n1271 , n1257 , n1270 , n1243 );
nand ( n1272 , n1269 , n1271 );
nor ( n1273 , n1264 , n1272 );
nand ( n1274 , n1250 , n1273 );
nand ( n1275 , n1230 , n1105 , n1047 );
not ( n1276 , n1275 );
not ( n1277 , n1237 );
not ( n1278 , n1277 );
and ( n1279 , n1276 , n1278 );
and ( n1280 , n149 , n1229 );
and ( n1281 , n1280 , n1247 );
and ( n1282 , n1281 , n1257 );
nor ( n1283 , n1279 , n1282 );
nand ( n1284 , n1047 , n1253 );
and ( n1285 , n1239 , n1280 );
nand ( n1286 , n1257 , n1285 , n1243 );
and ( n1287 , n1284 , n1286 );
nand ( n1288 , n1230 , n1239 , n1047 );
not ( n1289 , n1288 );
not ( n1290 , n1243 );
not ( n1291 , n1290 );
and ( n1292 , n1289 , n1291 );
and ( n1293 , n1001 , n1236 );
not ( n1294 , n1293 );
nor ( n1295 , n1234 , n1294 );
and ( n1296 , n1295 , n1257 );
nor ( n1297 , n1292 , n1296 );
and ( n1298 , n1283 , n1287 , n1297 );
nor ( n1299 , n1298 , n754 );
nor ( n1300 , n1274 , n1299 );
not ( n1301 , n754 );
nor ( n1302 , n35 , n31 , n1267 );
nand ( n1303 , n1301 , n1302 , n1247 );
not ( n1304 , n754 );
not ( n1305 , n1260 );
not ( n1306 , n1239 );
not ( n1307 , n1001 );
nor ( n1308 , n1305 , n1306 , n1307 );
nand ( n1309 , n1304 , n1257 , n1308 );
and ( n1310 , n1303 , n1309 );
nand ( n1311 , n1300 , n1310 );
nand ( n1312 , n1226 , n1311 );
nand ( n1313 , n140 , n1312 );
and ( n1314 , n20 , n1134 );
not ( n1315 , n1314 );
not ( n1316 , n724 );
nor ( n1317 , n1315 , n1316 );
and ( n1318 , n1313 , n1317 );
nor ( n1319 , n1315 , n295 );
not ( n1320 , n1129 );
and ( n1321 , n821 , n744 );
nand ( n1322 , n1302 , n1321 , n683 );
not ( n1323 , n675 );
nand ( n1324 , n1323 , n1308 , n683 );
nand ( n1325 , n1322 , n1324 );
not ( n1326 , n1325 );
nand ( n1327 , n1268 , n1321 , n1323 );
not ( n1328 , n678 );
not ( n1329 , n1328 );
nand ( n1330 , n1323 , n1270 , n1329 );
nand ( n1331 , n1327 , n1330 );
not ( n1332 , n1331 );
not ( n1333 , n822 );
and ( n1334 , n1095 , n1333 );
and ( n1335 , n1323 , n1334 , n1235 );
and ( n1336 , n1255 , n1323 );
nor ( n1337 , n1335 , n1336 );
buf ( n1338 , n1333 );
nand ( n1339 , n1260 , n1003 , n1338 );
and ( n1340 , n1242 , n678 );
and ( n1341 , n1245 , n1321 );
nor ( n1342 , n1340 , n1341 );
and ( n1343 , n1232 , n1339 , n1342 );
nand ( n1344 , n1332 , n1337 , n1343 );
not ( n1345 , n683 );
buf ( n1346 , n658 );
nor ( n1347 , n1346 , n1307 );
nand ( n1348 , n1233 , n1347 );
or ( n1349 , n1348 , n675 );
or ( n1350 , n1328 , n1288 );
nand ( n1351 , n1349 , n1350 );
nand ( n1352 , n1285 , n678 );
or ( n1353 , n675 , n1352 );
nand ( n1354 , n1353 , n1284 );
nand ( n1355 , n1280 , n1321 );
or ( n1356 , n675 , n1355 );
or ( n1357 , n1275 , n1346 );
nand ( n1358 , n1356 , n1357 );
nor ( n1359 , n1351 , n1354 , n1358 );
nor ( n1360 , n1345 , n1359 );
nor ( n1361 , n1344 , n1360 );
nand ( n1362 , n1326 , n1361 );
nand ( n1363 , n1320 , n1362 );
nand ( n1364 , n140 , n1363 );
and ( n1365 , n1319 , n1364 );
nor ( n1366 , n1318 , n1365 );
and ( n1367 , n1149 , n1224 , n1366 );
not ( n1368 , n18 );
not ( n1369 , n20 );
and ( n1370 , n1368 , n1369 );
not ( n1371 , n1370 );
nand ( n1372 , n16 , n19 );
not ( n1373 , n1372 );
and ( n1374 , n17 , n15 , n1373 );
not ( n1375 , n1374 );
nor ( n1376 , n1371 , n1375 );
not ( n1377 , n32 );
not ( n1378 , n134 );
nor ( n1379 , n25 , n1378 );
or ( n1380 , n1377 , n1379 );
not ( n1381 , n32 );
nor ( n1382 , n1381 , n26 );
not ( n1383 , n1382 );
nand ( n1384 , n1380 , n1383 );
not ( n1385 , n218 );
nand ( n1386 , n1384 , n153 , n1385 );
and ( n1387 , n32 , n26 , n234 );
and ( n1388 , n151 , n353 , n1387 );
nor ( n1389 , n1388 , n277 );
not ( n1390 , n266 );
nand ( n1391 , n355 , n1390 );
not ( n1392 , n1391 );
nand ( n1393 , n1392 , n575 );
and ( n1394 , n1386 , n1389 , n1393 );
or ( n1395 , n573 , n1394 );
nand ( n1396 , n1395 , n140 );
and ( n1397 , n1376 , n1396 );
not ( n1398 , n705 );
not ( n1399 , n17 );
nand ( n1400 , n22 , n1399 );
nand ( n1401 , n1398 , n1400 );
nand ( n1402 , n16 , n1401 );
nor ( n1403 , n1315 , n1402 );
nand ( n1404 , n19 , n1370 );
not ( n1405 , n18 );
and ( n1406 , n20 , n1405 );
or ( n1407 , n16 , n19 );
nand ( n1408 , n1372 , n1407 );
nand ( n1409 , n1406 , n1408 );
and ( n1410 , n1404 , n1409 );
not ( n1411 , n1401 );
nor ( n1412 , n1410 , n1411 );
nor ( n1413 , n1397 , n1403 , n1412 );
not ( n1414 , n18 );
nand ( n1415 , n1414 , n908 );
nor ( n1416 , n16 , n1415 );
nand ( n1417 , n1416 , n1401 );
nand ( n1418 , n20 , n781 );
nor ( n1419 , n18 , n1418 );
and ( n1420 , n1384 , n153 , n944 );
or ( n1421 , n945 , n1391 );
nand ( n1422 , n1421 , n1389 );
nor ( n1423 , n1420 , n1422 );
not ( n1424 , n1423 );
and ( n1425 , n525 , n1424 );
nor ( n1426 , n1425 , n139 );
not ( n1427 , n1426 );
and ( n1428 , n1419 , n1427 );
nor ( n1429 , n18 , n1411 );
and ( n1430 , n453 , n1429 );
nor ( n1431 , n1428 , n1430 );
nor ( n1432 , n18 , n523 );
not ( n1433 , n1130 );
not ( n1434 , n558 );
nand ( n1435 , n32 , n1053 );
nand ( n1436 , n209 , n1078 );
not ( n1437 , n1436 );
not ( n1438 , n1437 );
nand ( n1439 , n1435 , n1098 , n1001 , n1438 );
nor ( n1440 , n1434 , n1439 , n547 );
and ( n1441 , n548 , n1440 );
not ( n1442 , n1025 );
nand ( n1443 , n32 , n1442 );
nand ( n1444 , n1443 , n1160 , n1052 , n1438 );
buf ( n1445 , n541 );
not ( n1446 , n1445 );
and ( n1447 , n1028 , n1436 );
not ( n1448 , n1158 );
nand ( n1449 , n1052 , n1446 , n1447 , n1448 );
nand ( n1450 , n1444 , n1449 );
not ( n1451 , n547 );
and ( n1452 , n1450 , n1451 );
nor ( n1453 , n1441 , n1452 );
nand ( n1454 , n32 , n35 );
nor ( n1455 , n1454 , n1307 );
and ( n1456 , n1170 , n1447 , n1455 );
buf ( n1457 , n1445 );
and ( n1458 , n35 , n998 , n1051 );
and ( n1459 , n1458 , n1436 );
and ( n1460 , n1459 , n1098 , n409 );
not ( n1461 , n1027 );
and ( n1462 , n1435 , n1461 , n1458 , n1436 );
nor ( n1463 , n1460 , n1462 );
or ( n1464 , n1457 , n1463 );
not ( n1465 , n1437 );
not ( n1466 , n1065 );
nor ( n1467 , n1454 , n1053 , n1307 );
and ( n1468 , n1465 , n1466 , n1467 );
nor ( n1469 , n1468 , n411 );
nand ( n1470 , n1464 , n1469 );
nor ( n1471 , n1456 , n1470 );
not ( n1472 , n559 );
not ( n1473 , n1447 );
nor ( n1474 , n1169 , n1473 , n1457 );
not ( n1475 , n35 );
nor ( n1476 , n1475 , n23 );
and ( n1477 , n998 , n1476 );
nand ( n1478 , n1472 , n1474 , n1477 );
nand ( n1479 , n1453 , n1471 , n1478 );
not ( n1480 , n559 );
buf ( n1481 , n534 );
buf ( n1482 , n1481 );
and ( n1483 , n1158 , n1482 );
not ( n1484 , n540 );
nor ( n1485 , n1483 , n1484 );
not ( n1486 , n1012 );
nor ( n1487 , n31 , n1008 , n1486 );
not ( n1488 , n23 );
and ( n1489 , n1487 , n1488 , n1436 );
and ( n1490 , n1485 , n1451 , n1489 );
nand ( n1491 , n1443 , n1098 , n1477 , n1438 );
not ( n1492 , n1491 );
nor ( n1493 , n1490 , n1492 );
not ( n1494 , n1493 );
and ( n1495 , n1480 , n1494 );
nand ( n1496 , n1160 , n543 );
not ( n1497 , n1496 );
and ( n1498 , n1095 , n1438 );
not ( n1499 , n546 );
not ( n1500 , n1499 );
nand ( n1501 , n1497 , n1498 , n1500 );
buf ( n1502 , n532 );
buf ( n1503 , n1502 );
or ( n1504 , n1501 , n1503 , n1169 );
not ( n1505 , n1008 );
not ( n1506 , n23 );
and ( n1507 , n1436 , n1505 , n1506 );
not ( n1508 , n1065 );
not ( n1509 , n32 );
nor ( n1510 , n1509 , n31 );
and ( n1511 , n1507 , n1508 , n1510 );
nand ( n1512 , n1451 , n1511 , n1485 );
nand ( n1513 , n1504 , n1512 );
nor ( n1514 , n1495 , n1513 );
not ( n1515 , n1457 );
and ( n1516 , n1515 , n1447 , n558 );
nand ( n1517 , n1516 , n1451 , n153 , n1170 );
nand ( n1518 , n1001 , n1465 );
nor ( n1519 , n1496 , n1518 , n1499 );
nor ( n1520 , n1502 , n1158 );
and ( n1521 , n1519 , n1520 );
nand ( n1522 , n35 , n998 , n1066 , n1507 );
not ( n1523 , n1522 );
and ( n1524 , n1523 , n1485 );
nor ( n1525 , n1521 , n1524 );
not ( n1526 , n1525 );
not ( n1527 , n559 );
and ( n1528 , n1526 , n1527 );
and ( n1529 , n1438 , n1105 , n1477 );
and ( n1530 , n1529 , n1159 );
and ( n1531 , n1530 , n548 , n1103 , n558 );
nor ( n1532 , n1528 , n1531 );
nand ( n1533 , n1514 , n1517 , n1532 );
nor ( n1534 , n1479 , n1533 );
not ( n1535 , n1534 );
not ( n1536 , n1535 );
or ( n1537 , n1433 , n1536 );
nand ( n1538 , n1537 , n140 );
and ( n1539 , n1432 , n1538 );
not ( n1540 , n284 );
not ( n1541 , n20 );
nand ( n1542 , n1541 , n296 );
nor ( n1543 , n1540 , n1542 );
nor ( n1544 , n1539 , n1543 );
and ( n1545 , n1413 , n1417 , n1431 , n1544 );
not ( n1546 , n14 );
nor ( n1547 , n1546 , n20 );
not ( n1548 , n1547 );
nand ( n1549 , n18 , n430 );
nor ( n1550 , n1548 , n1549 );
not ( n1551 , n368 );
and ( n1552 , n1550 , n1551 );
not ( n1553 , n20 );
not ( n1554 , n294 );
nand ( n1555 , n1554 , n724 );
nor ( n1556 , n1553 , n1555 );
and ( n1557 , n1556 , n758 );
nor ( n1558 , n1552 , n1557 );
nor ( n1559 , n20 , n1555 );
and ( n1560 , n1559 , n510 );
nor ( n1561 , n14 , n20 );
not ( n1562 , n1549 );
nand ( n1563 , n1561 , n1562 );
nor ( n1564 , n1563 , n421 );
nor ( n1565 , n1560 , n1564 );
and ( n1566 , n1558 , n1565 );
not ( n1567 , n778 );
nand ( n1568 , n18 , n522 );
or ( n1569 , n1567 , n1568 );
not ( n1570 , n772 );
not ( n1571 , n591 );
nand ( n1572 , n18 , n1571 );
or ( n1573 , n1570 , n1572 );
nand ( n1574 , n1569 , n1573 );
nand ( n1575 , n18 , n908 );
not ( n1576 , n1575 );
not ( n1577 , n16 );
nand ( n1578 , n1577 , n1401 );
not ( n1579 , n1578 );
and ( n1580 , n1576 , n1579 );
nand ( n1581 , n19 , n309 );
and ( n1582 , n18 , n20 );
nand ( n1583 , n1582 , n1408 );
and ( n1584 , n1581 , n1583 );
nor ( n1585 , n1584 , n1411 );
nor ( n1586 , n1580 , n1585 );
not ( n1587 , n18 );
not ( n1588 , n20 );
nand ( n1589 , n1588 , n1374 );
nor ( n1590 , n1587 , n1589 );
and ( n1591 , n1590 , n784 );
nor ( n1592 , n971 , n1575 );
and ( n1593 , n1592 , n950 );
nor ( n1594 , n1591 , n1593 );
not ( n1595 , n18 );
nor ( n1596 , n1595 , n841 );
not ( n1597 , n16 );
not ( n1598 , n20 );
or ( n1599 , n1598 , n294 );
nor ( n1600 , n1597 , n1599 );
or ( n1601 , n1596 , n1600 );
nand ( n1602 , n1601 , n1401 );
not ( n1603 , n825 );
not ( n1604 , n1603 );
not ( n1605 , n831 );
and ( n1606 , n1604 , n1605 );
and ( n1607 , n796 , n805 );
nor ( n1608 , n1606 , n1607 );
nand ( n1609 , n870 , n1608 );
and ( n1610 , n1406 , n1609 );
not ( n1611 , n1141 );
nand ( n1612 , n1547 , n1611 );
not ( n1613 , n1612 );
not ( n1614 , n363 );
or ( n1615 , n943 , n1614 );
nand ( n1616 , n1615 , n140 );
and ( n1617 , n1613 , n1616 );
nor ( n1618 , n1610 , n1617 );
nand ( n1619 , n1586 , n1594 , n1602 , n1618 );
nor ( n1620 , n1574 , n1619 );
nor ( n1621 , n1575 , n521 );
and ( n1622 , n1621 , n906 );
nor ( n1623 , n1575 , n632 );
and ( n1624 , n1623 , n940 );
nor ( n1625 , n1622 , n1624 );
and ( n1626 , n872 , n1582 );
and ( n1627 , n20 , n296 );
and ( n1628 , n1627 , n688 );
nor ( n1629 , n1626 , n1628 );
and ( n1630 , n1620 , n1625 , n1629 );
not ( n1631 , n900 );
and ( n1632 , n206 , n1078 );
nor ( n1633 , n1632 , n1011 );
not ( n1634 , n1633 );
nor ( n1635 , n23 , n1634 );
and ( n1636 , n35 , n998 , n1635 );
not ( n1637 , n886 );
nor ( n1638 , n1637 , n798 );
nand ( n1639 , n1631 , n1636 , n1638 );
buf ( n1640 , n893 );
nand ( n1641 , n896 , n1640 );
buf ( n1642 , n894 );
not ( n1643 , n1642 );
nor ( n1644 , n1641 , n889 , n1643 );
not ( n1645 , n557 );
not ( n1646 , n1645 );
not ( n1647 , n1646 );
not ( n1648 , n1634 );
buf ( n1649 , n1648 );
not ( n1650 , n1505 );
not ( n1651 , n1650 );
and ( n1652 , n1649 , n1651 , n1001 );
nand ( n1653 , n1644 , n898 , n1647 , n1652 );
and ( n1654 , n1639 , n1653 );
not ( n1655 , n901 );
not ( n1656 , n1649 );
not ( n1657 , n1656 );
nand ( n1658 , n1657 , n1640 , n1642 );
nand ( n1659 , n896 , n1293 );
or ( n1660 , n1658 , n1659 );
nand ( n1661 , n1649 , n1651 , n1477 );
not ( n1662 , n888 );
or ( n1663 , n1661 , n1662 );
nand ( n1664 , n1660 , n1663 );
not ( n1665 , n1664 );
or ( n1666 , n1655 , n1665 );
nand ( n1667 , n1642 , n896 , n1640 );
and ( n1668 , n151 , n1648 );
nand ( n1669 , n1668 , n1638 );
or ( n1670 , n1667 , n1669 );
not ( n1671 , n1104 );
and ( n1672 , n1648 , n1671 , n1477 );
nand ( n1673 , n1672 , n1237 );
nand ( n1674 , n1670 , n1673 );
nand ( n1675 , n901 , n1674 );
nand ( n1676 , n1666 , n1675 );
not ( n1677 , n1676 );
and ( n1678 , n1443 , n1633 );
nand ( n1679 , n1477 , n1678 );
not ( n1680 , n1679 );
not ( n1681 , n896 );
not ( n1682 , n1650 );
nand ( n1683 , n1649 , n151 , n1682 );
nor ( n1684 , n1681 , n1683 );
not ( n1685 , n1662 );
nand ( n1686 , n1684 , n1685 , n1640 , n1642 );
not ( n1687 , n1686 );
or ( n1688 , n1680 , n1687 );
nand ( n1689 , n1688 , n901 );
nand ( n1690 , n1677 , n1689 );
not ( n1691 , n1467 );
not ( n1692 , n1648 );
or ( n1693 , n1691 , n1692 );
not ( n1694 , n277 );
nand ( n1695 , n1693 , n1694 );
not ( n1696 , n1695 );
nand ( n1697 , n1649 , n1455 , n1237 );
nand ( n1698 , n1458 , n1633 );
not ( n1699 , n1698 );
and ( n1700 , n1699 , n1638 );
nor ( n1701 , n1008 , n1698 );
not ( n1702 , n1701 );
nor ( n1703 , n1702 , n1662 );
nor ( n1704 , n1700 , n1703 );
nand ( n1705 , n1696 , n1697 , n1704 );
and ( n1706 , n32 , n998 , n1635 );
nand ( n1707 , n1706 , n1638 );
nand ( n1708 , n1642 , n896 , n1640 );
or ( n1709 , n1707 , n1708 );
nand ( n1710 , n1052 , n1678 );
nor ( n1711 , n1681 , n1710 );
nand ( n1712 , n1711 , n1640 , n1642 );
nand ( n1713 , n1709 , n1712 );
nor ( n1714 , n1705 , n1713 );
and ( n1715 , n896 , n1262 );
not ( n1716 , n1656 );
nand ( n1717 , n1715 , n1716 , n1640 , n1642 );
and ( n1718 , n1648 , n1505 , n1052 );
and ( n1719 , n896 , n1718 );
nand ( n1720 , n1719 , n1685 , n1640 , n1642 );
and ( n1721 , n1717 , n1720 );
nand ( n1722 , n1714 , n1721 );
nor ( n1723 , n1690 , n1722 );
nand ( n1724 , n1654 , n1723 );
not ( n1725 , n1225 );
and ( n1726 , n1724 , n1725 );
nor ( n1727 , n1726 , n139 );
buf ( n1728 , n1727 );
not ( n1729 , n1728 );
not ( n1730 , n1415 );
nand ( n1731 , n1729 , n1730 , n520 );
not ( n1732 , n1226 );
and ( n1733 , n608 , n1489 );
not ( n1734 , n600 );
nand ( n1735 , n1733 , n1734 , n602 , n596 );
nand ( n1736 , n1491 , n1735 );
and ( n1737 , n618 , n1736 );
nand ( n1738 , n1511 , n1734 , n596 );
not ( n1739 , n608 );
not ( n1740 , n602 );
or ( n1741 , n1738 , n1739 , n1740 );
nor ( n1742 , n1740 , n1067 );
nand ( n1743 , n1742 , n1498 , n596 );
nand ( n1744 , n608 , n1116 );
or ( n1745 , n1743 , n1744 );
nand ( n1746 , n1741 , n1745 );
nor ( n1747 , n1737 , n1746 );
not ( n1748 , n1518 );
nand ( n1749 , n1748 , n596 , n1068 , n602 );
nand ( n1750 , n608 , n1042 );
or ( n1751 , n1749 , n1750 );
not ( n1752 , n1734 );
or ( n1753 , n1522 , n1752 );
nand ( n1754 , n1751 , n1753 );
and ( n1755 , n618 , n1754 );
and ( n1756 , n615 , n1042 , n1160 , n1645 );
nand ( n1757 , n1756 , n1529 , n611 );
and ( n1758 , n596 , n608 , n602 );
and ( n1759 , n1447 , n1124 );
nor ( n1760 , n612 , n600 );
nand ( n1761 , n1758 , n1759 , n616 , n1760 );
nand ( n1762 , n1757 , n1761 );
nor ( n1763 , n1755 , n1762 );
and ( n1764 , n1747 , n1763 );
not ( n1765 , n617 );
not ( n1766 , n1752 );
and ( n1767 , n1766 , n1447 , n1017 );
nand ( n1768 , n1765 , n1767 , n1477 );
and ( n1769 , n1455 , n1447 , n1018 );
and ( n1770 , n1459 , n1098 , n1115 );
nor ( n1771 , n1770 , n1462 );
or ( n1772 , n1752 , n1771 );
nand ( n1773 , n1772 , n1469 );
nor ( n1774 , n1769 , n1773 );
nand ( n1775 , n608 , n602 , n615 , n596 );
nor ( n1776 , n1775 , n1646 , n1439 );
and ( n1777 , n611 , n1776 );
nand ( n1778 , n1052 , n1734 , n1447 , n1016 );
nand ( n1779 , n1444 , n1778 );
and ( n1780 , n1779 , n1758 );
nor ( n1781 , n1777 , n1780 );
and ( n1782 , n1768 , n1774 , n1781 );
nand ( n1783 , n1764 , n1782 );
not ( n1784 , n1783 );
or ( n1785 , n1732 , n1784 );
nand ( n1786 , n1785 , n140 );
nor ( n1787 , n18 , n591 );
and ( n1788 , n1786 , n1787 );
not ( n1789 , n1226 );
and ( n1790 , n918 , n925 , n928 );
nand ( n1791 , n1716 , n1334 , n1790 );
nand ( n1792 , n886 , n823 );
not ( n1793 , n1792 );
nand ( n1794 , n1706 , n1793 , n1790 );
nand ( n1795 , n1791 , n1794 );
not ( n1796 , n1795 );
not ( n1797 , n931 );
nor ( n1798 , n1797 , n929 );
nand ( n1799 , n930 , n1798 , n1647 , n1652 );
not ( n1800 , n929 );
not ( n1801 , n1710 );
and ( n1802 , n1800 , n1801 );
nor ( n1803 , n1802 , n1695 );
and ( n1804 , n1648 , n1455 , n1333 );
or ( n1805 , n1698 , n1792 );
not ( n1806 , n924 );
nand ( n1807 , n1701 , n1806 );
nand ( n1808 , n1805 , n1807 );
nor ( n1809 , n1804 , n1808 );
buf ( n1810 , n1806 );
nand ( n1811 , n1790 , n1718 , n1810 );
and ( n1812 , n1803 , n1809 , n1811 );
and ( n1813 , n1796 , n1799 , n1812 );
not ( n1814 , n932 );
not ( n1815 , n1810 );
or ( n1816 , n1815 , n1683 , n929 );
nand ( n1817 , n1816 , n1679 );
nand ( n1818 , n1814 , n1817 );
not ( n1819 , n932 );
nand ( n1820 , n1636 , n1793 , n1819 );
or ( n1821 , n1661 , n1815 );
nand ( n1822 , n1790 , n1347 , n1716 );
nand ( n1823 , n1821 , n1822 );
not ( n1824 , n1672 );
not ( n1825 , n1338 );
or ( n1826 , n1824 , n1825 );
nand ( n1827 , n1790 , n1793 , n1668 );
nand ( n1828 , n1826 , n1827 );
or ( n1829 , n1823 , n1828 );
nand ( n1830 , n1829 , n1814 );
nand ( n1831 , n1813 , n1818 , n1820 , n1830 );
not ( n1832 , n1831 );
not ( n1833 , n1832 );
not ( n1834 , n1833 );
or ( n1835 , n1789 , n1834 );
nand ( n1836 , n1835 , n140 );
nor ( n1837 , n1415 , n632 );
and ( n1838 , n1836 , n1837 );
nor ( n1839 , n1788 , n1838 );
and ( n1840 , n1566 , n1630 , n1731 , n1839 );
nand ( n1841 , n1367 , n1545 , n1840 );
not ( n1842 , n1841 );
not ( n1843 , n1842 );
and ( n1844 , n996 , n1843 );
not ( n1845 , n11 );
not ( n1846 , n13 );
nor ( n1847 , n1846 , n12 );
not ( n1848 , n1847 );
and ( n1849 , n1845 , n1848 );
nand ( n1850 , n1841 , n1849 );
nor ( n1851 , n11 , n12 );
and ( n1852 , n13 , n1851 );
or ( n1853 , n1407 , n1411 );
not ( n1854 , n103 );
nand ( n1855 , n1854 , n428 );
nand ( n1856 , n1853 , n1855 );
and ( n1857 , n1406 , n1856 );
not ( n1858 , n1730 );
not ( n1859 , n1722 );
nand ( n1860 , n1654 , n1859 , n1689 , n1677 );
not ( n1861 , n1860 );
or ( n1862 , n521 , n1861 );
nand ( n1863 , n1831 , n590 );
not ( n1864 , n102 );
not ( n1865 , n1864 );
not ( n1866 , n1865 );
not ( n1867 , n1866 );
not ( n1868 , n1867 );
not ( n1869 , n1868 );
not ( n1870 , n1869 );
not ( n1871 , n16 );
not ( n1872 , n448 );
nand ( n1873 , n1871 , n1872 );
or ( n1874 , n1870 , n1873 );
nand ( n1875 , n1874 , n1578 );
not ( n1876 , n1875 );
nand ( n1877 , n1862 , n1863 , n1876 );
not ( n1878 , n1877 );
or ( n1879 , n1858 , n1878 );
not ( n1880 , n583 );
or ( n1881 , n1534 , n1880 );
not ( n1882 , n1394 );
nand ( n1883 , n1374 , n1882 );
nand ( n1884 , n1881 , n1883 );
not ( n1885 , n1884 );
not ( n1886 , n1783 );
not ( n1887 , n1886 );
not ( n1888 , n764 );
not ( n1889 , n1888 );
and ( n1890 , n1887 , n1889 );
buf ( n1891 , n448 );
not ( n1892 , n1891 );
nand ( n1893 , n19 , n1892 );
or ( n1894 , n1870 , n1893 );
not ( n1895 , n19 );
nor ( n1896 , n1411 , n1895 );
not ( n1897 , n1896 );
nand ( n1898 , n1894 , n1897 );
nor ( n1899 , n1890 , n1898 );
nand ( n1900 , n1885 , n1899 );
not ( n1901 , n1900 );
or ( n1902 , n1901 , n1371 );
nand ( n1903 , n1879 , n1902 );
nor ( n1904 , n1857 , n1903 );
not ( n1905 , n1218 );
and ( n1906 , n1223 , n1905 );
and ( n1907 , n1137 , n1128 );
not ( n1908 , n20 );
nor ( n1909 , n1908 , n1222 );
not ( n1910 , n1909 );
not ( n1911 , n1311 );
or ( n1912 , n1910 , n1911 );
nand ( n1913 , n20 , n1136 );
not ( n1914 , n1362 );
buf ( n1915 , n1914 );
or ( n1916 , n1913 , n1915 );
nand ( n1917 , n1912 , n1916 );
nor ( n1918 , n1906 , n1907 , n1917 );
and ( n1919 , n20 , n1373 );
not ( n1920 , n1919 );
nor ( n1921 , n18 , n1920 );
and ( n1922 , n1921 , n1401 );
not ( n1923 , n1870 );
nor ( n1924 , n18 , n963 );
and ( n1925 , n1923 , n1924 );
nor ( n1926 , n1922 , n1925 );
not ( n1927 , n18 );
not ( n1928 , n22 );
nand ( n1929 , n23 , n428 );
or ( n1930 , n1928 , n20 , n1929 );
or ( n1931 , n16 , n841 );
or ( n1932 , n1931 , n1411 );
nand ( n1933 , n1930 , n1932 );
and ( n1934 , n1927 , n1933 );
or ( n1935 , n1143 , n1145 );
buf ( n1936 , n830 );
not ( n1937 , n1936 );
not ( n1938 , n1937 );
nand ( n1939 , n20 , n1938 );
nor ( n1940 , n18 , n1939 );
not ( n1941 , n1940 );
buf ( n1942 , n1603 );
not ( n1943 , n1942 );
buf ( n1944 , n1943 );
not ( n1945 , n1944 );
or ( n1946 , n1941 , n1945 );
nand ( n1947 , n20 , n1142 );
not ( n1948 , n1947 );
not ( n1949 , n805 );
not ( n1950 , n1949 );
and ( n1951 , n1948 , n1950 );
and ( n1952 , n1613 , n363 );
nor ( n1953 , n1951 , n1952 );
nand ( n1954 , n1935 , n1946 , n1953 );
not ( n1955 , n1419 );
not ( n1956 , n1424 );
or ( n1957 , n1955 , n1956 );
nor ( n1958 , n20 , n1135 );
or ( n1959 , n1314 , n1958 );
buf ( n1960 , n972 );
or ( n1961 , n1870 , n1960 );
nand ( n1962 , n1961 , n1402 );
nand ( n1963 , n1959 , n1962 );
nand ( n1964 , n1957 , n1963 );
nor ( n1965 , n1934 , n1954 , n1964 );
nand ( n1966 , n1904 , n1918 , n1926 , n1965 );
nand ( n1967 , n1852 , n1966 );
not ( n1968 , n1962 );
not ( n1969 , n1968 );
not ( n1970 , n20 );
not ( n1971 , n1852 );
nor ( n1972 , n294 , n1971 );
nand ( n1973 , n1969 , n1970 , n1972 );
not ( n1974 , n18 );
nor ( n1975 , n1974 , n1920 );
and ( n1976 , n1845 , n1847 );
and ( n1977 , n1975 , n1976 , n1401 );
and ( n1978 , n1592 , n1923 , n1852 );
nor ( n1979 , n1977 , n1978 );
not ( n1980 , n12 );
and ( n1981 , n13 , n1845 );
and ( n1982 , n18 , n1980 , n1981 );
and ( n1983 , n1982 , n1933 );
not ( n1984 , n1582 );
nor ( n1985 , n1984 , n1971 );
and ( n1986 , n1985 , n1856 );
nor ( n1987 , n1983 , n1986 );
nand ( n1988 , n1979 , n1987 );
nand ( n1989 , n18 , n942 );
or ( n1990 , n1971 , n1989 );
or ( n1991 , n1990 , n948 );
nand ( n1992 , n20 , n1972 );
or ( n1993 , n1992 , n1968 );
not ( n1994 , n1561 );
not ( n1995 , n431 );
not ( n1996 , n1995 );
nand ( n1997 , n1996 , n1982 );
nor ( n1998 , n1994 , n1997 );
not ( n1999 , n858 );
and ( n2000 , n1998 , n1999 );
not ( n2001 , n14 );
nand ( n2002 , n1582 , n431 );
nor ( n2003 , n2001 , n2002 );
and ( n2004 , n1852 , n2003 );
not ( n2005 , n827 );
and ( n2006 , n2004 , n2005 );
nor ( n2007 , n2000 , n2006 );
nand ( n2008 , n1991 , n1993 , n2007 );
nor ( n2009 , n20 , n294 );
and ( n2010 , n2009 , n1852 );
nand ( n2011 , n96 , n2010 );
not ( n2012 , n282 );
or ( n2013 , n2011 , n2012 );
nor ( n2014 , n1316 , n1599 , n1971 );
not ( n2015 , n2014 );
not ( n2016 , n756 );
or ( n2017 , n2015 , n2016 );
nor ( n2018 , n1548 , n1997 );
and ( n2019 , n2018 , n366 );
not ( n2020 , n14 );
not ( n2021 , n2002 );
nand ( n2022 , n2020 , n2021 );
nor ( n2023 , n1971 , n2022 );
and ( n2024 , n2023 , n808 );
nor ( n2025 , n2019 , n2024 );
nand ( n2026 , n2013 , n2017 , n2025 );
nor ( n2027 , n1988 , n2008 , n2026 );
and ( n2028 , n724 , n2010 );
and ( n2029 , n2028 , n506 );
nor ( n2030 , n1971 , n1599 , n295 );
and ( n2031 , n2030 , n686 );
nor ( n2032 , n2029 , n2031 );
nor ( n2033 , n308 , n1971 );
and ( n2034 , n764 , n621 );
nor ( n2035 , n2034 , n1898 );
and ( n2036 , n583 , n564 );
and ( n2037 , n1374 , n579 );
nor ( n2038 , n2036 , n2037 );
nand ( n2039 , n2035 , n2038 );
and ( n2040 , n2033 , n2039 );
nor ( n2041 , n1575 , n1971 );
not ( n2042 , n520 );
not ( n2043 , n904 );
or ( n2044 , n2042 , n2043 );
and ( n2045 , n590 , n936 );
nor ( n2046 , n2045 , n1875 );
nand ( n2047 , n2044 , n2046 );
and ( n2048 , n2041 , n2047 );
nor ( n2049 , n2040 , n2048 );
and ( n2050 , n2027 , n2032 , n2049 );
nand ( n2051 , n1850 , n1967 , n1973 , n2050 );
not ( n2052 , n2 );
and ( n2053 , n2051 , n2052 );
nor ( n2054 , n1844 , n2053 );
nand ( n2055 , n787 , n637 , n442 );
not ( n2056 , n289 );
not ( n2057 , n1836 );
or ( n2058 , n2057 , n913 );
or ( n2059 , n963 , n1426 );
nand ( n2060 , n2058 , n2059 );
nor ( n2061 , n1728 , n910 );
nor ( n2062 , n2060 , n2061 );
or ( n2063 , n2056 , n2062 );
not ( n2064 , n90 );
not ( n2065 , n450 );
and ( n2066 , n16 , n642 );
not ( n2067 , n2066 );
nor ( n2068 , n2065 , n2067 );
nand ( n2069 , n2064 , n2068 );
not ( n2070 , n2069 );
buf ( n2071 , n1313 );
and ( n2072 , n2070 , n2071 );
not ( n2073 , n20 );
nor ( n2074 , n2073 , n90 );
and ( n2075 , n2074 , n1609 );
nor ( n2076 , n2072 , n2075 );
nor ( n2077 , n41 , n868 );
nand ( n2078 , n812 , n1608 );
nand ( n2079 , n2077 , n2078 );
not ( n2080 , n633 );
not ( n2081 , n975 );
not ( n2082 , n2081 );
and ( n2083 , n2080 , n2082 );
not ( n2084 , n1724 );
or ( n2085 , n2084 , n955 );
or ( n2086 , n961 , n1832 );
nand ( n2087 , n2085 , n2086 );
nor ( n2088 , n2083 , n2087 );
and ( n2089 , n965 , n1424 );
and ( n2090 , n909 , n811 );
nor ( n2091 , n2089 , n2090 );
nand ( n2092 , n2088 , n2091 );
and ( n2093 , n2056 , n2092 );
and ( n2094 , n20 , n99 );
and ( n2095 , n2094 , n1364 );
nor ( n2096 , n2093 , n2095 );
nand ( n2097 , n2063 , n2076 , n2079 , n2096 );
nand ( n2098 , n286 , n2068 );
and ( n2099 , n300 , n1312 );
or ( n2100 , n2098 , n2099 );
not ( n2101 , n20 );
nand ( n2102 , n90 , n97 );
nor ( n2103 , n2101 , n2102 );
not ( n2104 , n2103 );
and ( n2105 , n300 , n1363 );
or ( n2106 , n2104 , n2105 );
not ( n2107 , n20 );
not ( n2108 , n306 );
or ( n2109 , n2107 , n2108 );
nand ( n2110 , n2109 , n912 );
and ( n2111 , n2110 , n334 );
nor ( n2112 , n692 , n330 );
or ( n2113 , n318 , n2112 );
not ( n2114 , n14 );
nand ( n2115 , n2113 , n2114 );
not ( n2116 , n2115 );
and ( n2117 , n2066 , n2116 );
nor ( n2118 , n2111 , n2117 );
nand ( n2119 , n2100 , n2106 , n2118 );
or ( n2120 , n2097 , n2119 );
nor ( n2121 , n18 , n81 );
nand ( n2122 , n2120 , n2121 );
not ( n2123 , n795 );
and ( n2124 , n2123 , n1147 );
buf ( n2125 , n1938 );
not ( n2126 , n2125 );
not ( n2127 , n2126 );
buf ( n2128 , n2127 );
and ( n2129 , n2128 , n1616 );
nor ( n2130 , n2124 , n2129 );
not ( n2131 , n2130 );
nand ( n2132 , n853 , n2131 );
nand ( n2133 , n300 , n1220 );
and ( n2134 , n838 , n2133 );
not ( n2135 , n796 );
not ( n2136 , n415 );
or ( n2137 , n2135 , n2136 );
not ( n2138 , n831 );
not ( n2139 , n1614 );
and ( n2140 , n2138 , n2139 );
nor ( n2141 , n2140 , n813 );
nand ( n2142 , n2137 , n2141 );
and ( n2143 , n856 , n2142 );
nor ( n2144 , n2134 , n2143 );
and ( n2145 , n790 , n1221 );
and ( n2146 , n1132 , n848 );
nor ( n2147 , n2145 , n2146 );
and ( n2148 , n2132 , n2144 , n2147 );
not ( n2149 , n851 );
not ( n2150 , n40 );
not ( n2151 , n2150 );
not ( n2152 , n1535 );
not ( n2153 , n2152 );
and ( n2154 , n2153 , n527 );
buf ( n2155 , n1783 );
and ( n2156 , n592 , n2155 );
nor ( n2157 , n2154 , n2156 );
not ( n2158 , n634 );
and ( n2159 , n574 , n1882 );
nor ( n2160 , n2159 , n586 );
and ( n2161 , n2157 , n2158 , n2160 );
not ( n2162 , n2161 );
and ( n2163 , n2151 , n2162 );
not ( n2164 , n40 );
not ( n2165 , n2164 );
not ( n2166 , n584 );
not ( n2167 , n1538 );
or ( n2168 , n2166 , n2167 );
and ( n2169 , n1786 , n1571 );
and ( n2170 , n570 , n1396 );
nor ( n2171 , n2169 , n2170 );
nand ( n2172 , n2168 , n2171 );
not ( n2173 , n2172 );
or ( n2174 , n2165 , n2173 );
nand ( n2175 , n300 , n1131 );
nand ( n2176 , n844 , n2175 );
nand ( n2177 , n2174 , n2176 );
nor ( n2178 , n2163 , n2177 );
nand ( n2179 , n2148 , n2149 , n2178 );
not ( n2180 , n18 );
not ( n2181 , n988 );
nand ( n2182 , n2180 , n2181 );
not ( n2183 , n2182 );
nand ( n2184 , n2179 , n2183 );
and ( n2185 , n2055 , n2122 , n2184 );
not ( n2186 , n454 );
not ( n2187 , n442 );
or ( n2188 , n2115 , n2186 , n2187 );
not ( n2189 , n628 );
not ( n2190 , n2189 );
not ( n2191 , n2190 );
not ( n2192 , n2191 );
not ( n2193 , n2192 );
not ( n2194 , n2193 );
not ( n2195 , n2194 );
not ( n2196 , n2195 );
or ( n2197 , n2196 , n333 , n2187 );
nand ( n2198 , n2188 , n2197 );
nand ( n2199 , n445 , n853 );
or ( n2200 , n863 , n2199 , n2187 );
not ( n2201 , n2118 );
not ( n2202 , n2074 );
not ( n2203 , n872 );
or ( n2204 , n2202 , n2203 );
or ( n2205 , n2098 , n876 );
nand ( n2206 , n2204 , n2205 );
nor ( n2207 , n2201 , n2206 );
not ( n2208 , n833 );
nand ( n2209 , n2208 , n2077 );
and ( n2210 , n2103 , n719 );
and ( n2211 , n2094 , n688 );
nor ( n2212 , n2210 , n2211 );
and ( n2213 , n289 , n953 );
not ( n2214 , n288 );
not ( n2215 , n910 );
not ( n2216 , n905 );
and ( n2217 , n2215 , n2216 );
nor ( n2218 , n2217 , n977 );
or ( n2219 , n2214 , n2218 );
or ( n2220 , n2069 , n759 );
nand ( n2221 , n2219 , n2220 );
nor ( n2222 , n2213 , n2221 );
and ( n2223 , n2207 , n2209 , n2212 , n2222 );
or ( n2224 , n2223 , n2187 );
nand ( n2225 , n2200 , n2224 );
nor ( n2226 , n2198 , n2225 );
not ( n2227 , n14 );
or ( n2228 , n2227 , n447 );
not ( n2229 , n2228 );
nand ( n2230 , n2229 , n454 );
nor ( n2231 , n40 , n2230 );
and ( n2232 , n445 , n2231 );
and ( n2233 , n2232 , n2175 );
nand ( n2234 , n14 , n16 );
not ( n2235 , n2234 );
or ( n2236 , n2235 , n841 );
nand ( n2237 , n2236 , n2192 );
and ( n2238 , n2237 , n334 );
not ( n2239 , n16 );
not ( n2240 , n19 );
nand ( n2241 , n2240 , n1547 );
or ( n2242 , n2239 , n2241 );
not ( n2243 , n2242 );
nand ( n2244 , n14 , n17 );
not ( n2245 , n2244 );
nand ( n2246 , n92 , n2245 );
or ( n2247 , n2246 , n330 );
nand ( n2248 , n2247 , n319 );
and ( n2249 , n2243 , n2248 );
nor ( n2250 , n2233 , n2238 , n2249 );
buf ( n2251 , n2172 );
and ( n2252 , n291 , n2251 );
or ( n2253 , n2161 , n291 );
not ( n2254 , n2133 );
not ( n2255 , n789 );
nand ( n2256 , n288 , n2255 );
or ( n2257 , n2254 , n2256 );
nand ( n2258 , n2253 , n2257 );
nor ( n2259 , n2252 , n2258 );
and ( n2260 , n440 , n2131 );
nand ( n2261 , n2245 , n454 );
not ( n2262 , n331 );
or ( n2263 , n2261 , n2262 );
not ( n2264 , n2199 );
nand ( n2265 , n2264 , n2142 );
nand ( n2266 , n2263 , n2265 );
nor ( n2267 , n2260 , n2266 );
nor ( n2268 , n288 , n789 );
and ( n2269 , n2268 , n1221 );
nor ( n2270 , n286 , n2230 );
and ( n2271 , n2270 , n1132 );
nor ( n2272 , n2269 , n2271 );
and ( n2273 , n2267 , n2272 );
and ( n2274 , n2250 , n2259 , n2273 );
not ( n2275 , n2121 );
nor ( n2276 , n2274 , n2275 );
and ( n2277 , n40 , n2092 );
or ( n2278 , n2062 , n40 );
or ( n2279 , n717 , n2105 );
nand ( n2280 , n2278 , n2279 );
nor ( n2281 , n2277 , n2280 );
not ( n2282 , n714 );
not ( n2283 , n794 );
nand ( n2284 , n2283 , n2078 );
not ( n2285 , n2099 );
and ( n2286 , n875 , n2285 );
and ( n2287 , n869 , n1609 );
nor ( n2288 , n2286 , n2287 );
and ( n2289 , n726 , n2071 );
and ( n2290 , n648 , n1364 );
nor ( n2291 , n2289 , n2290 );
and ( n2292 , n2284 , n2288 , n2291 );
and ( n2293 , n2281 , n2282 , n2292 );
nor ( n2294 , n2293 , n2182 );
nor ( n2295 , n2276 , n2294 );
nand ( n2296 , n2054 , n2185 , n2226 , n2295 );
or ( n2297 , n991 , n2296 );
not ( n2298 , n3 );
not ( n2299 , n5 );
and ( n2300 , n2298 , n2299 );
and ( n2301 , n1 , n2300 );
nand ( n2302 , n2297 , n2301 );
not ( n2303 , n42 );
nor ( n2304 , n2303 , n725 );
and ( n2305 , n2304 , n756 );
or ( n2306 , n42 , n795 );
not ( n2307 , n40 );
and ( n2308 , n41 , n2307 );
not ( n2309 , n2308 );
not ( n2310 , n2309 );
not ( n2311 , n2310 );
not ( n2312 , n2311 );
not ( n2313 , n2312 );
not ( n2314 , n26 );
nor ( n2315 , n2314 , n25 );
not ( n2316 , n2315 );
buf ( n2317 , n2316 );
not ( n2318 , n2317 );
not ( n2319 , n224 );
or ( n2320 , n2318 , n2319 );
nor ( n2321 , n148 , n227 );
nand ( n2322 , n2320 , n2321 );
not ( n2323 , n2322 );
or ( n2324 , n22 , n2323 );
and ( n2325 , n2313 , n2324 );
not ( n2326 , n2313 );
and ( n2327 , n275 , n2322 );
nand ( n2328 , n299 , n2327 );
and ( n2329 , n2326 , n2328 );
nor ( n2330 , n2325 , n2329 );
or ( n2331 , n2306 , n2330 );
not ( n2332 , n1407 );
not ( n2333 , n22 );
not ( n2334 , n2312 );
and ( n2335 , n2333 , n2334 );
not ( n2336 , n2312 );
not ( n2337 , n314 );
or ( n2338 , n2336 , n2337 );
not ( n2339 , n17 );
nand ( n2340 , n2338 , n2339 );
nor ( n2341 , n2335 , n2340 );
not ( n2342 , n2341 );
not ( n2343 , n14 );
nand ( n2344 , n2343 , n17 );
not ( n2345 , n2344 );
not ( n2346 , n2345 );
not ( n2347 , n2346 );
not ( n2348 , n2347 );
not ( n2349 , n2348 );
not ( n2350 , n2311 );
and ( n2351 , n2350 , n326 );
and ( n2352 , n2311 , n328 );
nor ( n2353 , n2351 , n2352 );
nor ( n2354 , n15 , n2353 );
nand ( n2355 , n2349 , n2354 );
nand ( n2356 , n2342 , n2355 );
and ( n2357 , n2332 , n2356 );
not ( n2358 , n2334 );
not ( n2359 , n2358 );
or ( n2360 , n2359 , n299 );
not ( n2361 , n2334 );
or ( n2362 , n1868 , n2361 );
nand ( n2363 , n2360 , n2362 );
not ( n2364 , n2363 );
nor ( n2365 , n2303 , n2364 );
and ( n2366 , n2123 , n2365 );
nor ( n2367 , n2357 , n2366 );
nand ( n2368 , n2331 , n2367 );
and ( n2369 , n20 , n2368 );
nor ( n2370 , n42 , n2330 );
or ( n2371 , n2365 , n2370 );
and ( n2372 , n590 , n2371 );
not ( n2373 , n16 );
or ( n2374 , n2246 , n2353 );
not ( n2375 , n2341 );
nand ( n2376 , n2374 , n2375 );
and ( n2377 , n2373 , n2376 );
nor ( n2378 , n2372 , n2377 );
nor ( n2379 , n912 , n2378 );
nor ( n2380 , n2305 , n2369 , n2379 );
not ( n2381 , n20 );
nor ( n2382 , n2381 , n14 );
not ( n2383 , n19 );
or ( n2384 , n2383 , n16 );
not ( n2385 , n2384 );
nand ( n2386 , n2382 , n2385 );
nand ( n2387 , n14 , n20 );
nor ( n2388 , n19 , n2387 );
and ( n2389 , n16 , n2388 );
not ( n2390 , n2388 );
or ( n2391 , n16 , n2390 );
not ( n2392 , n2391 );
nor ( n2393 , n2389 , n2392 );
nand ( n2394 , n2386 , n2393 );
not ( n2395 , n448 );
nand ( n2396 , n2303 , n2395 );
or ( n2397 , n2396 , n2330 );
nor ( n2398 , n2303 , n448 );
and ( n2399 , n2398 , n2363 );
nor ( n2400 , n692 , n2353 );
nor ( n2401 , n2399 , n2400 );
nand ( n2402 , n2397 , n2401 );
and ( n2403 , n2394 , n2402 );
not ( n2404 , n2371 );
nor ( n2405 , n963 , n2404 );
nor ( n2406 , n2403 , n2405 );
not ( n2407 , n970 );
nand ( n2408 , n42 , n2407 );
nor ( n2409 , n912 , n2408 );
nand ( n2410 , n2409 , n966 );
and ( n2411 , n2354 , n17 );
nor ( n2412 , n2411 , n2341 );
not ( n2413 , n2412 );
nand ( n2414 , n1919 , n2413 );
nand ( n2415 , n2380 , n2406 , n2410 , n2414 );
not ( n2416 , n431 );
nor ( n2417 , n1994 , n2416 );
and ( n2418 , n42 , n2417 );
not ( n2419 , n2418 );
buf ( n2420 , n1999 );
not ( n2421 , n2420 );
or ( n2422 , n2419 , n2421 );
and ( n2423 , n724 , n2371 );
and ( n2424 , n16 , n2356 );
nor ( n2425 , n2423 , n2424 );
or ( n2426 , n841 , n2425 );
and ( n2427 , n2243 , n2402 );
and ( n2428 , n570 , n2371 );
nor ( n2429 , n2427 , n2428 );
nand ( n2430 , n2422 , n2426 , n2429 );
nand ( n2431 , n2398 , n2392 );
or ( n2432 , n2431 , n827 );
not ( n2433 , n646 );
not ( n2434 , n2433 );
not ( n2435 , n2434 );
not ( n2436 , n2435 );
not ( n2437 , n2436 );
not ( n2438 , n2437 );
not ( n2439 , n2438 );
not ( n2440 , n2439 );
not ( n2441 , n2440 );
or ( n2442 , n2441 , n2425 );
not ( n2443 , n2398 );
not ( n2444 , n16 );
not ( n2445 , n2241 );
nand ( n2446 , n2444 , n2445 );
nor ( n2447 , n2443 , n2446 );
and ( n2448 , n2447 , n366 );
not ( n2449 , n20 );
or ( n2450 , n2303 , n795 );
nor ( n2451 , n2449 , n2450 );
and ( n2452 , n2451 , n808 );
nor ( n2453 , n2448 , n2452 );
nand ( n2454 , n2432 , n2442 , n2453 );
nor ( n2455 , n2415 , n2430 , n2454 );
not ( n2456 , n16 );
not ( n2457 , n623 );
and ( n2458 , n2456 , n2457 );
and ( n2459 , n2458 , n2356 );
not ( n2460 , n20 );
and ( n2461 , n42 , n2460 );
nand ( n2462 , n2461 , n781 );
not ( n2463 , n2462 );
nand ( n2464 , n2463 , n579 );
not ( n2465 , n20 );
and ( n2466 , n2465 , n2368 );
nand ( n2467 , n2385 , n1547 );
nand ( n2468 , n2467 , n2446 );
and ( n2469 , n2468 , n2402 );
nor ( n2470 , n2466 , n2469 );
nand ( n2471 , n2464 , n2470 );
not ( n2472 , n16 );
nor ( n2473 , n2472 , n2194 , n2412 );
not ( n2474 , n2473 );
nor ( n2475 , n2443 , n2467 );
nand ( n2476 , n2475 , n621 );
nand ( n2477 , n522 , n2371 );
nor ( n2478 , n2443 , n2242 );
nand ( n2479 , n2478 , n282 );
nand ( n2480 , n2474 , n2476 , n2477 , n2479 );
nor ( n2481 , n2459 , n2471 , n2480 );
nor ( n2482 , n2443 , n2386 );
buf ( n2483 , n958 );
not ( n2484 , n2483 );
and ( n2485 , n2482 , n2484 );
not ( n2486 , n20 );
nor ( n2487 , n2486 , n2303 );
nand ( n2488 , n19 , n2487 );
nor ( n2489 , n2488 , n632 );
not ( n2490 , n960 );
and ( n2491 , n2489 , n2490 );
nor ( n2492 , n2485 , n2491 );
nand ( n2493 , n2398 , n2389 );
not ( n2494 , n2493 );
not ( n2495 , n686 );
not ( n2496 , n2495 );
and ( n2497 , n2494 , n2496 );
or ( n2498 , n2303 , n521 );
or ( n2499 , n565 , n2190 , n2498 );
not ( n2500 , n506 );
nand ( n2501 , n42 , n724 );
or ( n2502 , n2500 , n841 , n2501 );
nand ( n2503 , n2499 , n2502 );
nor ( n2504 , n2497 , n2503 );
nand ( n2505 , n2455 , n2481 , n2492 , n2504 );
not ( n2506 , n1 );
and ( n2507 , n2506 , n2298 );
and ( n2508 , n2 , n2507 );
not ( n2509 , n2508 );
nor ( n2510 , n5 , n2509 );
nand ( n2511 , n2505 , n1982 , n2510 );
not ( n2512 , n2152 );
buf ( n2513 , n2512 );
buf ( n2514 , n2513 );
and ( n2515 , n2385 , n1561 );
not ( n2516 , n18 );
and ( n2517 , n2516 , n1980 , n1981 );
nand ( n2518 , n2517 , n2510 );
nor ( n2519 , n2443 , n2518 );
and ( n2520 , n2514 , n2515 , n2519 );
not ( n2521 , n2414 );
nor ( n2522 , n2521 , n2405 );
not ( n2523 , n2522 );
and ( n2524 , n96 , n2371 );
and ( n2525 , n16 , n2376 );
nor ( n2526 , n2524 , n2525 );
or ( n2527 , n2441 , n2526 );
not ( n2528 , n19 );
nand ( n2529 , n2528 , n2382 );
nor ( n2530 , n16 , n2529 );
nand ( n2531 , n805 , n2398 , n2530 );
nand ( n2532 , n2527 , n2531 );
not ( n2533 , n20 );
buf ( n2534 , n2128 );
and ( n2535 , n2534 , n2370 );
and ( n2536 , n2332 , n2376 );
nand ( n2537 , n14 , n42 );
nor ( n2538 , n2537 , n429 );
and ( n2539 , n2538 , n2363 );
nor ( n2540 , n2535 , n2536 , n2539 );
or ( n2541 , n2533 , n2540 );
not ( n2542 , n972 );
not ( n2543 , n2488 );
and ( n2544 , n2542 , n2543 );
nand ( n2545 , n2544 , n1424 );
nand ( n2546 , n2541 , n2545 );
nor ( n2547 , n2523 , n2532 , n2546 , n2379 );
not ( n2548 , n16 );
nor ( n2549 , n2548 , n2529 );
and ( n2550 , n1311 , n2398 , n2549 );
nand ( n2551 , n20 , n2538 );
not ( n2552 , n1944 );
or ( n2553 , n2551 , n2552 );
nand ( n2554 , n42 , n590 );
or ( n2555 , n1832 , n912 , n2554 );
nand ( n2556 , n2553 , n2555 );
nor ( n2557 , n2550 , n2556 );
and ( n2558 , n2530 , n2402 );
nor ( n2559 , n2303 , n647 );
not ( n2560 , n1915 );
nand ( n2561 , n2559 , n2560 );
nand ( n2562 , n2482 , n1724 );
nand ( n2563 , n2561 , n2562 );
not ( n2564 , n2549 );
and ( n2565 , n2386 , n2564 );
not ( n2566 , n2402 );
nor ( n2567 , n2565 , n2566 );
nor ( n2568 , n2558 , n2563 , n2567 );
and ( n2569 , n2547 , n2557 , n2568 );
nor ( n2570 , n2569 , n2518 );
nor ( n2571 , n2520 , n2570 );
and ( n2572 , n2302 , n2511 , n2571 );
not ( n2573 , n2230 );
not ( n2574 , n2358 );
not ( n2575 , n2574 );
not ( n2576 , n2575 );
not ( n2577 , n2576 );
not ( n2578 , n2 );
not ( n2579 , n1982 );
nor ( n2580 , n2578 , n2579 );
not ( n2581 , n2580 );
nor ( n2582 , n2577 , n2581 );
nand ( n2583 , n2573 , n2582 );
not ( n2584 , n2583 );
not ( n2585 , n1540 );
and ( n2586 , n2584 , n2585 );
not ( n2587 , n301 );
nand ( n2588 , n41 , n2580 , n2231 );
nor ( n2589 , n2587 , n2588 );
nor ( n2590 , n2586 , n2589 );
not ( n2591 , n2590 );
nand ( n2592 , n454 , n2580 );
or ( n2593 , n2341 , n2400 );
nand ( n2594 , n2593 , n14 );
or ( n2595 , n2592 , n2594 );
nand ( n2596 , n2193 , n2580 );
or ( n2597 , n2596 , n2412 );
nand ( n2598 , n2595 , n2597 );
not ( n2599 , n19 );
nand ( n2600 , n2599 , n2234 );
not ( n2601 , n20 );
nand ( n2602 , n2601 , n1982 );
not ( n2603 , n2602 );
nand ( n2604 , n2 , n2603 );
or ( n2605 , n2412 , n2600 , n2604 );
not ( n2606 , n20 );
not ( n2607 , n2575 );
nand ( n2608 , n2606 , n2607 );
nor ( n2609 , n2608 , n2581 );
not ( n2610 , n2609 );
not ( n2611 , n439 );
or ( n2612 , n2610 , n2611 );
nand ( n2613 , n2605 , n2612 );
not ( n2614 , n19 );
and ( n2615 , n2614 , n724 );
not ( n2616 , n2615 );
nor ( n2617 , n20 , n2616 );
and ( n2618 , n2617 , n2582 );
not ( n2619 , n2618 );
not ( n2620 , n510 );
or ( n2621 , n2619 , n2620 );
not ( n2622 , n20 );
not ( n2623 , n2576 );
nand ( n2624 , n2623 , n2615 );
not ( n2625 , n2624 );
nand ( n2626 , n2622 , n2580 , n2625 , n508 );
nand ( n2627 , n2621 , n2626 );
nor ( n2628 , n2591 , n2598 , n2613 , n2627 );
or ( n2629 , n2228 , n2067 );
nor ( n2630 , n2575 , n2629 );
and ( n2631 , n2630 , n1364 );
not ( n2632 , n20 );
nor ( n2633 , n2632 , n2575 );
and ( n2634 , n2633 , n1609 );
nor ( n2635 , n2631 , n2634 );
not ( n2636 , n2623 );
not ( n2637 , n2636 );
or ( n2638 , n2637 , n2062 );
or ( n2639 , n2576 , n725 );
or ( n2640 , n2639 , n2099 );
nand ( n2641 , n2637 , n2092 );
nand ( n2642 , n2638 , n2640 , n2641 );
not ( n2643 , n2642 );
and ( n2644 , n2635 , n2643 );
nor ( n2645 , n445 , n868 );
nand ( n2646 , n2645 , n2078 );
or ( n2647 , n2067 , n2594 );
not ( n2648 , n20 );
nor ( n2649 , n2648 , n2600 );
or ( n2650 , n908 , n2649 );
nand ( n2651 , n2650 , n2413 );
nand ( n2652 , n2647 , n2651 );
nor ( n2653 , n40 , n2629 );
nand ( n2654 , n41 , n2653 );
or ( n2655 , n2654 , n2105 );
or ( n2656 , n2577 , n725 );
not ( n2657 , n2071 );
or ( n2658 , n2656 , n2657 );
nand ( n2659 , n2655 , n2658 );
nor ( n2660 , n2652 , n2659 );
and ( n2661 , n2644 , n2646 , n2660 );
nand ( n2662 , n2 , n2517 );
nor ( n2663 , n2661 , n2662 );
nor ( n2664 , n2576 , n843 );
and ( n2665 , n2664 , n2175 );
nand ( n2666 , n41 , n456 );
nor ( n2667 , n2666 , n2254 );
or ( n2668 , n2608 , n2130 );
or ( n2669 , n2186 , n2355 );
not ( n2670 , n853 );
nor ( n2671 , n445 , n2670 );
nand ( n2672 , n2671 , n2142 );
nand ( n2673 , n2668 , n2669 , n2672 );
nor ( n2674 , n2665 , n2667 , n2673 );
nor ( n2675 , n2577 , n455 );
and ( n2676 , n2675 , n1221 );
nor ( n2677 , n19 , n1994 );
nand ( n2678 , n16 , n2677 );
not ( n2679 , n2678 );
and ( n2680 , n2679 , n2356 );
nand ( n2681 , n305 , n453 );
and ( n2682 , n2194 , n2681 );
nor ( n2683 , n2682 , n2412 );
nor ( n2684 , n2676 , n2680 , n2683 );
not ( n2685 , n2637 );
and ( n2686 , n2685 , n2251 );
or ( n2687 , n2161 , n2685 );
nand ( n2688 , n2576 , n842 );
not ( n2689 , n1132 );
or ( n2690 , n2688 , n2689 );
nand ( n2691 , n2687 , n2690 );
nor ( n2692 , n2686 , n2691 );
and ( n2693 , n2674 , n2684 , n2692 );
nor ( n2694 , n2693 , n2662 );
nor ( n2695 , n2663 , n2694 );
not ( n2696 , n2 );
nor ( n2697 , n2696 , n1976 );
and ( n2698 , n2697 , n1841 );
not ( n2699 , n2636 );
nand ( n2700 , n2699 , n2580 );
not ( n2701 , n2700 );
and ( n2702 , n2701 , n636 );
nor ( n2703 , n2698 , n2702 );
not ( n2704 , n2645 );
or ( n2705 , n2704 , n833 );
not ( n2706 , n2633 );
not ( n2707 , n872 );
or ( n2708 , n2706 , n2707 );
or ( n2709 , n2654 , n720 );
nand ( n2710 , n2708 , n2709 );
nor ( n2711 , n2652 , n2710 );
and ( n2712 , n2636 , n953 );
or ( n2713 , n2639 , n876 );
or ( n2714 , n2656 , n759 );
nand ( n2715 , n2713 , n2714 );
not ( n2716 , n2630 );
not ( n2717 , n688 );
or ( n2718 , n2716 , n2717 );
not ( n2719 , n2623 );
or ( n2720 , n2719 , n2218 );
nand ( n2721 , n2718 , n2720 );
nor ( n2722 , n2712 , n2715 , n2721 );
nand ( n2723 , n2705 , n2711 , n2722 );
and ( n2724 , n2723 , n2580 );
and ( n2725 , n2582 , n787 );
and ( n2726 , n2671 , n2580 );
and ( n2727 , n2726 , n864 );
nor ( n2728 , n2724 , n2725 , n2727 );
and ( n2729 , n2695 , n2703 , n2728 );
and ( n2730 , n2628 , n2729 );
not ( n2731 , n2301 );
nor ( n2732 , n2730 , n2731 );
not ( n2733 , n2196 );
not ( n2734 , n2518 );
nand ( n2735 , n2733 , n2734 );
not ( n2736 , n2554 );
nand ( n2737 , n1783 , n2736 );
or ( n2738 , n2735 , n2737 );
nand ( n2739 , n1905 , n2679 , n2519 );
nand ( n2740 , n2738 , n2739 );
and ( n2741 , n2303 , n1400 , n704 );
nor ( n2742 , n2741 , n20 );
and ( n2743 , n2039 , n2742 , n18 );
nand ( n2744 , n15 , n42 );
or ( n2745 , n2744 , n2346 );
nor ( n2746 , n19 , n1371 );
nand ( n2747 , n16 , n2746 );
nor ( n2748 , n2745 , n2747 );
and ( n2749 , n1905 , n2748 );
nor ( n2750 , n2743 , n2749 );
not ( n2751 , n18 );
not ( n2752 , n2543 );
not ( n2753 , n2047 );
or ( n2754 , n2752 , n2753 );
nand ( n2755 , n2754 , n2410 );
not ( n2756 , n2755 );
or ( n2757 , n2751 , n2756 );
not ( n2758 , n19 );
and ( n2759 , n2758 , n17 , n588 );
nor ( n2760 , n2759 , n1996 );
nand ( n2761 , n2303 , n2324 );
or ( n2762 , n2760 , n2761 );
and ( n2763 , n306 , n1401 );
not ( n2764 , n19 );
nand ( n2765 , n2764 , n1867 );
nand ( n2766 , n42 , n2229 );
or ( n2767 , n2765 , n2766 );
or ( n2768 , n2303 , n1855 );
nand ( n2769 , n2767 , n2768 );
nor ( n2770 , n2763 , n2769 );
nand ( n2771 , n2762 , n2770 );
nand ( n2772 , n1370 , n2771 );
nand ( n2773 , n2757 , n2772 );
not ( n2774 , n2761 );
and ( n2775 , n2774 , n450 );
nand ( n2776 , n1867 , n2398 );
and ( n2777 , n2776 , n1411 );
nor ( n2778 , n2777 , n14 );
nor ( n2779 , n2775 , n2778 );
or ( n2780 , n2747 , n2779 );
buf ( n2781 , n1891 );
or ( n2782 , n2781 , n2761 );
nand ( n2783 , n2782 , n2777 );
not ( n2784 , n2783 );
or ( n2785 , n1575 , n2784 );
nand ( n2786 , n2780 , n2785 );
nor ( n2787 , n2773 , n2786 );
not ( n2788 , n18 );
nand ( n2789 , n42 , n97 );
or ( n2790 , n2789 , n2495 );
not ( n2791 , n2538 );
not ( n2792 , n2791 );
not ( n2793 , n827 );
and ( n2794 , n2792 , n2793 );
nor ( n2795 , n807 , n2450 );
nor ( n2796 , n2794 , n2795 );
nand ( n2797 , n2790 , n2796 );
and ( n2798 , n20 , n2797 );
not ( n2799 , n20 );
nor ( n2800 , n2616 , n2303 );
nand ( n2801 , n2800 , n506 );
not ( n2802 , n2450 );
and ( n2803 , n2802 , n419 );
and ( n2804 , n366 , n2538 );
nor ( n2805 , n2803 , n2804 );
nand ( n2806 , n2801 , n2805 );
and ( n2807 , n2799 , n2806 );
nor ( n2808 , n2798 , n2807 );
or ( n2809 , n2788 , n2808 );
not ( n2810 , n18 );
nand ( n2811 , n1900 , n2742 , n2810 );
and ( n2812 , n2750 , n2787 , n2809 , n2811 );
nand ( n2813 , n1877 , n2543 );
not ( n2814 , n16 );
or ( n2815 , n2814 , n19 );
not ( n2816 , n2815 );
not ( n2817 , n20 );
nor ( n2818 , n2817 , n2745 );
nand ( n2819 , n1311 , n2816 , n2818 );
and ( n2820 , n20 , n2771 );
and ( n2821 , n908 , n2783 );
nor ( n2822 , n2820 , n2821 );
nand ( n2823 , n2813 , n2819 , n2822 );
not ( n2824 , n2823 );
or ( n2825 , n1914 , n2789 );
and ( n2826 , n2802 , n805 );
not ( n2827 , n1942 );
and ( n2828 , n2538 , n2827 );
nor ( n2829 , n2826 , n2828 );
nand ( n2830 , n2825 , n2829 );
nand ( n2831 , n20 , n2830 );
and ( n2832 , n2545 , n2831 );
not ( n2833 , n2779 );
nand ( n2834 , n2066 , n2833 );
nand ( n2835 , n2824 , n2832 , n2834 );
not ( n2836 , n18 );
and ( n2837 , n2835 , n2836 );
not ( n2838 , n2766 );
and ( n2839 , n282 , n2838 );
not ( n2840 , n2777 );
and ( n2841 , n14 , n2840 );
nor ( n2842 , n2839 , n2841 );
nand ( n2843 , n2816 , n309 );
or ( n2844 , n2842 , n2843 );
not ( n2845 , n434 );
and ( n2846 , n309 , n2845 );
and ( n2847 , n450 , n1596 );
nor ( n2848 , n2846 , n2847 );
or ( n2849 , n2848 , n2761 );
or ( n2850 , n1145 , n2450 );
nand ( n2851 , n2538 , n363 );
nand ( n2852 , n2850 , n2851 );
and ( n2853 , n1370 , n2852 );
or ( n2854 , n1411 , n2600 );
or ( n2855 , n2765 , n2745 );
nand ( n2856 , n2854 , n2855 , n2768 );
and ( n2857 , n309 , n2856 );
nor ( n2858 , n2853 , n2857 );
not ( n2859 , n2858 );
not ( n2860 , n16 );
not ( n2861 , n19 );
nand ( n2862 , n2861 , n1582 );
nor ( n2863 , n2860 , n2862 );
not ( n2864 , n2863 );
or ( n2865 , n2016 , n2745 , n2864 );
nor ( n2866 , n308 , n2228 );
and ( n2867 , n2816 , n2866 );
nor ( n2868 , n20 , n1893 );
nor ( n2869 , n2867 , n2868 );
or ( n2870 , n2869 , n2761 );
nand ( n2871 , n2865 , n2870 );
nor ( n2872 , n2859 , n2871 );
nand ( n2873 , n2844 , n2849 , n2872 );
not ( n2874 , n2873 );
and ( n2875 , n1582 , n2771 );
and ( n2876 , n2863 , n2833 );
nor ( n2877 , n2875 , n2876 );
not ( n2878 , n19 );
and ( n2879 , n42 , n2878 );
nand ( n2880 , n2879 , n96 , n1370 , n1128 );
nand ( n2881 , n2874 , n2877 , n2880 );
nor ( n2882 , n2837 , n2881 );
nand ( n2883 , n2812 , n2882 );
buf ( n2884 , n2883 );
not ( n2885 , n1976 );
and ( n2886 , n2884 , n2885 , n2510 );
nor ( n2887 , n2732 , n2740 , n2886 );
not ( n2888 , n2300 );
nor ( n2889 , n1 , n2888 );
not ( n2890 , n2889 );
not ( n2891 , n1849 );
not ( n2892 , n2883 );
or ( n2893 , n2891 , n2892 );
not ( n2894 , n20 );
nor ( n2895 , n42 , n2579 );
nor ( n2896 , n22 , n23 );
nand ( n2897 , n21 , n24 );
not ( n2898 , n2897 );
nand ( n2899 , n24 , n136 );
nand ( n2900 , n2896 , n998 , n2898 , n2899 );
and ( n2901 , n106 , n2900 );
not ( n2902 , n2899 );
and ( n2903 , n21 , n2902 );
not ( n2904 , n2903 );
nand ( n2905 , n2904 , n621 );
nand ( n2906 , n2901 , n2905 );
and ( n2907 , n764 , n2906 );
nor ( n2908 , n2907 , n1896 );
or ( n2909 , n565 , n2903 );
nand ( n2910 , n2909 , n2901 );
and ( n2911 , n583 , n2910 );
or ( n2912 , n2903 , n578 );
nand ( n2913 , n2912 , n2901 );
and ( n2914 , n1374 , n2913 );
nor ( n2915 , n2911 , n2914 );
nand ( n2916 , n2908 , n2915 );
nand ( n2917 , n2894 , n2895 , n2916 );
nand ( n2918 , n2893 , n2917 );
not ( n2919 , n2517 );
nor ( n2920 , n42 , n912 );
not ( n2921 , n2920 );
nor ( n2922 , n1832 , n2903 );
not ( n2923 , n2901 );
nor ( n2924 , n2922 , n2923 );
or ( n2925 , n632 , n2924 );
not ( n2926 , n2904 );
not ( n2927 , n1724 );
or ( n2928 , n2926 , n2927 );
nand ( n2929 , n2928 , n2901 );
nand ( n2930 , n2929 , n520 );
nand ( n2931 , n2925 , n2930 , n1578 );
not ( n2932 , n2931 );
or ( n2933 , n2921 , n2932 );
nand ( n2934 , n2933 , n2819 );
nand ( n2935 , n1311 , n2904 );
nand ( n2936 , n2901 , n2935 );
or ( n2937 , n92 , n42 );
nor ( n2938 , n2348 , n2937 );
and ( n2939 , n2936 , n2066 , n2938 );
nor ( n2940 , n2934 , n2939 );
nand ( n2941 , n2904 , n1362 );
and ( n2942 , n2901 , n2941 );
or ( n2943 , n2942 , n98 );
nand ( n2944 , n435 , n2923 );
not ( n2945 , n1936 );
nor ( n2946 , n2945 , n2903 );
nand ( n2947 , n2946 , n1943 );
nor ( n2948 , n795 , n2903 );
nand ( n2949 , n2948 , n805 );
and ( n2950 , n2944 , n2947 , n2949 );
nand ( n2951 , n2943 , n2950 );
not ( n2952 , n2951 );
not ( n2953 , n20 );
nor ( n2954 , n2953 , n42 );
not ( n2955 , n2954 );
nor ( n2956 , n2952 , n2955 );
or ( n2957 , n912 , n2777 );
or ( n2958 , n2903 , n1423 );
nand ( n2959 , n2958 , n2901 );
nand ( n2960 , n2959 , n2954 , n781 );
nand ( n2961 , n2957 , n2831 , n2960 );
not ( n2962 , n20 );
or ( n2963 , n2962 , n2770 );
nand ( n2964 , n2066 , n2778 );
nand ( n2965 , n2963 , n2964 , n2813 );
nor ( n2966 , n2956 , n2961 , n2965 );
nand ( n2967 , n2940 , n2545 , n2966 );
not ( n2968 , n2967 );
or ( n2969 , n2919 , n2968 );
not ( n2970 , n1901 );
not ( n2971 , n2461 );
not ( n2972 , n2971 );
and ( n2973 , n2970 , n2972 );
nand ( n2974 , n1128 , n2904 );
and ( n2975 , n2901 , n2974 );
not ( n2976 , n2975 );
nor ( n2977 , n42 , n2228 );
and ( n2978 , n454 , n2977 );
and ( n2979 , n2976 , n2978 );
nor ( n2980 , n2973 , n2979 );
not ( n2981 , n2904 );
not ( n2982 , n1535 );
or ( n2983 , n2981 , n2982 );
nand ( n2984 , n2983 , n2901 );
and ( n2985 , n2984 , n583 );
or ( n2986 , n2903 , n1394 );
nand ( n2987 , n2986 , n2901 );
and ( n2988 , n1374 , n2987 );
nor ( n2989 , n2985 , n2988 );
not ( n2990 , n2904 );
not ( n2991 , n1783 );
or ( n2992 , n2990 , n2991 );
nand ( n2993 , n2992 , n2901 );
and ( n2994 , n764 , n2993 );
nor ( n2995 , n2994 , n1896 );
nand ( n2996 , n2989 , n2995 );
not ( n2997 , n20 );
and ( n2998 , n2997 , n2303 );
nand ( n2999 , n2996 , n2998 );
not ( n3000 , n20 );
not ( n3001 , n2856 );
not ( n3002 , n3001 );
and ( n3003 , n3000 , n3002 );
not ( n3004 , n2615 );
not ( n3005 , n2904 );
not ( n3006 , n1217 );
or ( n3007 , n3005 , n3006 );
nand ( n3008 , n3007 , n2901 );
not ( n3009 , n3008 );
or ( n3010 , n3004 , n3009 );
or ( n3011 , n2903 , n1145 );
nand ( n3012 , n3011 , n2901 );
and ( n3013 , n2123 , n3012 );
or ( n3014 , n2903 , n1614 );
nand ( n3015 , n3014 , n2901 );
and ( n3016 , n2128 , n3015 );
nor ( n3017 , n3013 , n3016 );
nand ( n3018 , n3010 , n3017 );
and ( n3019 , n3018 , n2998 );
nor ( n3020 , n3003 , n3019 );
nand ( n3021 , n2243 , n2840 );
not ( n3022 , n20 );
nand ( n3023 , n3022 , n2852 );
nand ( n3024 , n1128 , n454 , n2838 );
nor ( n3025 , n2303 , n789 );
nand ( n3026 , n3025 , n1219 );
and ( n3027 , n3021 , n3023 , n3024 , n3026 );
nand ( n3028 , n2980 , n2999 , n3020 , n3027 );
nand ( n3029 , n3028 , n2517 );
nand ( n3030 , n2969 , n3029 );
nor ( n3031 , n2918 , n3030 );
nand ( n3032 , n2904 , n282 );
nand ( n3033 , n2901 , n3032 );
not ( n3034 , n3033 );
nand ( n3035 , n2977 , n1982 );
or ( n3036 , n3034 , n2186 , n3035 );
or ( n3037 , n2842 , n2815 , n2602 );
nand ( n3038 , n3036 , n3037 );
or ( n3039 , n2579 , n2808 );
nand ( n3040 , n2904 , n506 );
and ( n3041 , n2901 , n3040 );
or ( n3042 , n2616 , n3041 );
not ( n3043 , n14 );
or ( n3044 , n2903 , n365 );
nand ( n3045 , n3044 , n2901 );
or ( n3046 , n3043 , n3045 );
or ( n3047 , n857 , n2903 );
nand ( n3048 , n3047 , n2901 );
or ( n3049 , n14 , n3048 );
not ( n3050 , n436 );
nand ( n3051 , n3046 , n3049 , n3050 );
nand ( n3052 , n3042 , n3051 );
nand ( n3053 , n3052 , n2998 , n1982 );
nand ( n3054 , n3039 , n3053 );
nor ( n3055 , n3038 , n3054 );
and ( n3056 , n20 , n2895 );
not ( n3057 , n97 );
nand ( n3058 , n2904 , n686 );
nand ( n3059 , n2901 , n3058 );
not ( n3060 , n3059 );
or ( n3061 , n3057 , n3060 );
nand ( n3062 , n2948 , n808 );
nand ( n3063 , n2946 , n2005 );
and ( n3064 , n3062 , n2944 , n3063 );
nand ( n3065 , n3061 , n3064 );
and ( n3066 , n3056 , n3065 );
and ( n3067 , n1982 , n2755 );
nor ( n3068 , n3066 , n3067 );
and ( n3069 , n20 , n1982 );
not ( n3070 , n3069 );
not ( n3071 , n3070 );
not ( n3072 , n2770 );
and ( n3073 , n3071 , n3072 );
nor ( n3074 , n912 , n2579 );
and ( n3075 , n3074 , n2840 );
nor ( n3076 , n3073 , n3075 );
nand ( n3077 , n2904 , n756 );
nand ( n3078 , n2901 , n3077 );
nand ( n3079 , n2066 , n1982 );
not ( n3080 , n3079 );
and ( n3081 , n3078 , n2938 , n3080 );
not ( n3082 , n2745 );
and ( n3083 , n756 , n3082 , n3080 );
nor ( n3084 , n3081 , n3083 );
and ( n3085 , n2039 , n2461 , n1982 );
and ( n3086 , n3069 , n2816 , n2778 );
nor ( n3087 , n3085 , n3086 );
not ( n3088 , n16 );
nand ( n3089 , n3088 , n908 );
not ( n3090 , n3089 );
not ( n3091 , n3090 );
not ( n3092 , n1401 );
or ( n3093 , n3091 , n3092 );
not ( n3094 , n942 );
or ( n3095 , n2903 , n948 );
nand ( n3096 , n3095 , n2901 );
not ( n3097 , n3096 );
or ( n3098 , n3094 , n3097 );
or ( n3099 , n956 , n2903 );
nand ( n3100 , n3099 , n2901 );
and ( n3101 , n909 , n3100 );
nand ( n3102 , n2904 , n936 );
and ( n3103 , n3102 , n2901 );
nor ( n3104 , n3103 , n913 );
nor ( n3105 , n3101 , n3104 );
nand ( n3106 , n3098 , n3105 );
not ( n3107 , n3106 );
nand ( n3108 , n3093 , n3107 );
and ( n3109 , n3108 , n2895 );
and ( n3110 , n2603 , n2856 );
nor ( n3111 , n3109 , n3110 );
and ( n3112 , n3076 , n3084 , n3087 , n3111 );
nand ( n3113 , n3031 , n3055 , n3068 , n3112 );
not ( n3114 , n2 );
and ( n3115 , n3113 , n3114 );
not ( n3116 , n2 );
and ( n3117 , n11 , n1980 );
nand ( n3118 , n3116 , n3117 );
not ( n3119 , n3118 );
not ( n3120 , n3119 );
nor ( n3121 , n13 , n18 );
not ( n3122 , n3121 );
nand ( n3123 , n2512 , n2398 , n2515 );
nor ( n3124 , n2303 , n295 );
nand ( n3125 , n1128 , n3124 );
nor ( n3126 , n3125 , n841 );
not ( n3127 , n3126 );
not ( n3128 , n2515 );
nand ( n3129 , n3128 , n2678 );
not ( n3130 , n89 );
and ( n3131 , n3130 , n2324 );
not ( n3132 , n3130 );
and ( n3133 , n3132 , n2328 );
nor ( n3134 , n3131 , n3133 );
or ( n3135 , n3134 , n2396 );
not ( n3136 , n2443 );
not ( n3137 , n299 );
and ( n3138 , n89 , n3137 );
and ( n3139 , n1865 , n88 );
nor ( n3140 , n3138 , n3139 );
not ( n3141 , n3140 );
and ( n3142 , n3136 , n3141 );
nor ( n3143 , n3142 , n2112 );
nand ( n3144 , n3135 , n3143 );
and ( n3145 , n3129 , n3144 );
not ( n3146 , n2446 );
and ( n3147 , n3146 , n3144 );
nor ( n3148 , n3145 , n3147 );
and ( n3149 , n3123 , n3127 , n3148 );
nor ( n3150 , n2443 , n2678 );
nand ( n3151 , n3150 , n1905 );
nand ( n3152 , n2418 , n415 );
or ( n3153 , n2192 , n2737 );
and ( n3154 , n3151 , n3152 , n3153 );
or ( n3155 , n3134 , n42 );
or ( n3156 , n2303 , n3140 );
nand ( n3157 , n3155 , n3156 );
not ( n3158 , n3157 );
not ( n3159 , n3158 );
and ( n3160 , n96 , n3159 );
and ( n3161 , n16 , n2248 );
nor ( n3162 , n3160 , n3161 );
or ( n3163 , n841 , n3162 );
not ( n3164 , n20 );
or ( n3165 , n2306 , n3134 );
and ( n3166 , n2347 , n331 );
nor ( n3167 , n3166 , n318 );
or ( n3168 , n1407 , n3167 );
or ( n3169 , n795 , n3156 );
nand ( n3170 , n3165 , n3168 , n3169 );
and ( n3171 , n3164 , n3170 );
nor ( n3172 , n2462 , n1394 );
nor ( n3173 , n3171 , n3172 );
nand ( n3174 , n3163 , n3173 );
not ( n3175 , n630 );
not ( n3176 , n3175 );
and ( n3177 , n3157 , n590 );
not ( n3178 , n16 );
and ( n3179 , n3178 , n2248 );
nor ( n3180 , n3177 , n3179 );
or ( n3181 , n3176 , n3180 );
not ( n3182 , n2447 );
or ( n3183 , n3182 , n1614 );
not ( n3184 , n16 );
not ( n3185 , n627 );
not ( n3186 , n3185 );
or ( n3187 , n3184 , n3186 , n333 );
not ( n3188 , n3157 );
or ( n3189 , n3188 , n571 );
nand ( n3190 , n3187 , n3189 );
not ( n3191 , n3190 );
nand ( n3192 , n3181 , n3183 , n3191 );
nor ( n3193 , n3174 , n3192 );
nand ( n3194 , n3149 , n3154 , n3193 );
not ( n3195 , n3194 );
or ( n3196 , n3122 , n3195 );
nor ( n3197 , n13 , n1984 );
nand ( n3198 , n3197 , n2795 );
nand ( n3199 , n3196 , n3198 );
not ( n3200 , n2545 );
or ( n3201 , n2493 , n1915 );
not ( n3202 , n20 );
not ( n3203 , n3170 );
or ( n3204 , n3202 , n3203 );
nand ( n3205 , n3201 , n3204 , n2555 );
nor ( n3206 , n3200 , n3205 );
and ( n3207 , n2394 , n3144 );
or ( n3208 , n1316 , n3158 );
not ( n3209 , n16 );
or ( n3210 , n3209 , n3167 );
nand ( n3211 , n3208 , n3210 );
and ( n3212 , n2436 , n3211 );
not ( n3213 , n3180 );
and ( n3214 , n908 , n3213 );
nor ( n3215 , n3212 , n3214 );
nand ( n3216 , n2304 , n1311 );
nand ( n3217 , n3215 , n2562 , n3216 );
or ( n3218 , n2431 , n2552 );
not ( n3219 , n3159 );
or ( n3220 , n963 , n3219 );
and ( n3221 , n2487 , n2123 );
and ( n3222 , n3221 , n805 );
and ( n3223 , n1919 , n334 );
nor ( n3224 , n3222 , n3223 );
nand ( n3225 , n3218 , n3220 , n3224 );
nor ( n3226 , n3207 , n3217 , n3225 );
and ( n3227 , n3206 , n3226 );
not ( n3228 , n3121 );
nor ( n3229 , n3227 , n3228 );
nor ( n3230 , n3199 , n3229 );
and ( n3231 , n3197 , n3170 );
nor ( n3232 , n305 , n13 , n2862 );
not ( n3233 , n3232 );
or ( n3234 , n2016 , n2443 , n3233 );
not ( n3235 , n13 );
nand ( n3236 , n18 , n3235 );
nor ( n3237 , n19 , n3236 );
nand ( n3238 , n20 , n3237 );
not ( n3239 , n3124 );
or ( n3240 , n2495 , n3238 , n3239 );
nand ( n3241 , n3234 , n3240 );
not ( n3242 , n1575 );
not ( n3243 , n3242 );
not ( n3244 , n13 );
not ( n3245 , n14 );
nor ( n3246 , n3245 , n16 );
nand ( n3247 , n3244 , n3246 );
nor ( n3248 , n3243 , n3247 , n960 , n2443 );
nor ( n3249 , n3231 , n3241 , n3248 );
not ( n3250 , n3236 );
not ( n3251 , n2467 );
or ( n3252 , n3251 , n2243 );
nand ( n3253 , n3252 , n3144 );
not ( n3254 , n2503 );
and ( n3255 , n2479 , n2476 , n3253 , n3254 );
not ( n3256 , n1931 );
and ( n3257 , n3256 , n2248 );
or ( n3258 , n521 , n3158 );
or ( n3259 , n16 , n3167 );
nand ( n3260 , n3258 , n3259 );
not ( n3261 , n3260 );
or ( n3262 , n3176 , n3261 );
not ( n3263 , n20 );
nand ( n3264 , n3263 , n1936 );
nor ( n3265 , n42 , n3264 );
not ( n3266 , n3134 );
and ( n3267 , n3265 , n3266 );
nor ( n3268 , n3267 , n3190 );
nand ( n3269 , n3262 , n3268 );
nand ( n3270 , n2461 , n2125 );
or ( n3271 , n3270 , n3140 );
nand ( n3272 , n3271 , n2464 );
nor ( n3273 , n3257 , n3269 , n3272 );
not ( n3274 , n16 );
nand ( n3275 , n3274 , n2677 );
nor ( n3276 , n2443 , n3275 );
and ( n3277 , n3276 , n2420 );
not ( n3278 , n3275 );
and ( n3279 , n3278 , n3144 );
nor ( n3280 , n3277 , n3279 );
not ( n3281 , n3270 );
and ( n3282 , n3281 , n366 );
and ( n3283 , n453 , n3211 );
nor ( n3284 , n3282 , n3283 );
nand ( n3285 , n3255 , n3273 , n3280 , n3284 );
and ( n3286 , n3250 , n3285 );
not ( n3287 , n13 );
nand ( n3288 , n3287 , n3242 );
nor ( n3289 , n2483 , n3288 , n2498 );
nor ( n3290 , n3286 , n3289 );
or ( n3291 , n3238 , n3162 );
not ( n3292 , n3288 );
and ( n3293 , n3246 , n3292 );
nor ( n3294 , n3293 , n3232 );
not ( n3295 , n3144 );
or ( n3296 , n3294 , n3295 );
not ( n3297 , n19 );
nand ( n3298 , n14 , n3297 );
nor ( n3299 , n16 , n3298 );
and ( n3300 , n3144 , n3197 , n3299 );
and ( n3301 , n3292 , n3260 );
nor ( n3302 , n3300 , n3301 );
nand ( n3303 , n3291 , n3296 , n3302 );
or ( n3304 , n3219 , n13 , n1989 );
not ( n3305 , n2544 );
or ( n3306 , n948 , n3236 , n3305 );
nand ( n3307 , n3304 , n3306 );
not ( n3308 , n3197 );
nand ( n3309 , n2398 , n3299 );
or ( n3310 , n827 , n3308 , n3309 );
not ( n3311 , n1975 );
or ( n3312 , n13 , n3311 , n333 );
nand ( n3313 , n3310 , n3312 );
nor ( n3314 , n3303 , n3307 , n3313 );
nand ( n3315 , n3230 , n3249 , n3290 , n3314 );
not ( n3316 , n3315 );
or ( n3317 , n3120 , n3316 );
not ( n3318 , n40 );
and ( n3319 , n3318 , n2324 );
not ( n3320 , n3318 );
and ( n3321 , n3320 , n2328 );
nor ( n3322 , n3319 , n3321 );
or ( n3323 , n3322 , n42 );
and ( n3324 , n40 , n3137 );
not ( n3325 , n40 );
and ( n3326 , n3325 , n1867 );
nor ( n3327 , n3324 , n3326 );
or ( n3328 , n2303 , n3327 );
nand ( n3329 , n3323 , n3328 );
nand ( n3330 , n782 , n3329 );
not ( n3331 , n1960 );
buf ( n3332 , n3331 );
and ( n3333 , n3332 , n3329 );
not ( n3334 , n713 );
and ( n3335 , n16 , n3334 );
nor ( n3336 , n3333 , n3335 );
nor ( n3337 , n841 , n3336 );
not ( n3338 , n3337 );
and ( n3339 , n433 , n3329 );
and ( n3340 , n2332 , n3334 );
nor ( n3341 , n3339 , n3340 );
nor ( n3342 , n20 , n3341 );
not ( n3343 , n3342 );
nand ( n3344 , n3330 , n3338 , n3343 , n3023 );
nor ( n3345 , n20 , n1372 );
not ( n3346 , n3345 );
nor ( n3347 , n3346 , n713 );
nor ( n3348 , n3344 , n3347 , n3172 );
nand ( n3349 , n42 , n583 );
nor ( n3350 , n20 , n3349 );
and ( n3351 , n3350 , n2513 );
not ( n3352 , n1873 );
and ( n3353 , n3352 , n3329 );
not ( n3354 , n16 );
and ( n3355 , n3354 , n3334 );
nor ( n3356 , n3353 , n3355 );
nor ( n3357 , n3176 , n3356 );
not ( n3358 , n3127 );
nor ( n3359 , n3351 , n3357 , n3358 );
nand ( n3360 , n3153 , n3026 , n3348 , n3359 );
nand ( n3361 , n2183 , n3360 );
nand ( n3362 , n3317 , n3361 );
nor ( n3363 , n3115 , n3362 );
not ( n3364 , n989 );
nor ( n3365 , n2439 , n3336 );
not ( n3366 , n3365 );
or ( n3367 , n3364 , n3366 );
not ( n3368 , n988 );
not ( n3369 , n3368 );
not ( n3370 , n3369 );
not ( n3371 , n3370 );
not ( n3372 , n3371 );
not ( n3373 , n3372 );
not ( n3374 , n3373 );
nand ( n3375 , n1582 , n3374 );
or ( n3376 , n3375 , n3341 );
nand ( n3377 , n3367 , n3376 );
not ( n3378 , n994 );
not ( n3379 , n2883 );
or ( n3380 , n3378 , n3379 );
not ( n3381 , n3356 );
not ( n3382 , n3373 );
not ( n3383 , n3382 );
not ( n3384 , n3383 );
nand ( n3385 , n3381 , n3242 , n3384 );
nand ( n3386 , n3380 , n3385 );
nor ( n3387 , n3377 , n3386 );
not ( n3388 , n20 );
or ( n3389 , n3388 , n3341 );
or ( n3390 , n1920 , n713 );
nand ( n3391 , n3389 , n3390 , n2545 );
not ( n3392 , n20 );
or ( n3393 , n3392 , n2829 );
or ( n3394 , n912 , n3356 );
not ( n3395 , n3329 );
or ( n3396 , n963 , n3395 );
nand ( n3397 , n3393 , n3394 , n3396 );
nor ( n3398 , n3391 , n3397 );
nor ( n3399 , n2488 , n521 );
not ( n3400 , n2084 );
and ( n3401 , n3399 , n3400 );
not ( n3402 , n3216 );
nor ( n3403 , n3401 , n3365 , n3402 );
nand ( n3404 , n3398 , n3403 , n2555 , n2561 );
and ( n3405 , n2183 , n3404 );
or ( n3406 , n20 , n2805 );
nand ( n3407 , n42 , n626 );
or ( n3408 , n1960 , n3407 );
or ( n3409 , n3408 , n578 );
not ( n3410 , n3347 );
nor ( n3411 , n3357 , n3337 , n3342 );
nand ( n3412 , n3410 , n3411 , n3330 );
nor ( n3413 , n2971 , n1888 );
not ( n3414 , n3413 );
not ( n3415 , n621 );
or ( n3416 , n3414 , n3415 );
nand ( n3417 , n42 , n842 );
or ( n3418 , n3417 , n2012 );
nand ( n3419 , n3416 , n3418 , n3254 );
nor ( n3420 , n3412 , n3419 );
nand ( n3421 , n3406 , n3409 , n3420 );
and ( n3422 , n3421 , n989 );
nor ( n3423 , n3405 , n3422 );
nand ( n3424 , n3242 , n3382 , n2736 , n2490 );
not ( n3425 , n1599 );
not ( n3426 , n2501 );
nand ( n3427 , n3425 , n3382 , n3426 , n756 );
nor ( n3428 , n3369 , n3239 );
nand ( n3429 , n686 , n3425 , n3428 );
not ( n3430 , n2498 );
nand ( n3431 , n3242 , n3382 , n3430 , n2484 );
nand ( n3432 , n3424 , n3427 , n3429 , n3431 );
not ( n3433 , n18 );
not ( n3434 , n3332 );
not ( n3435 , n3434 );
not ( n3436 , n3435 );
nor ( n3437 , n3433 , n3436 );
nand ( n3438 , n3437 , n3329 );
or ( n3439 , n3438 , n912 , n3383 );
not ( n3440 , n989 );
or ( n3441 , n948 , n3440 , n3305 );
nand ( n3442 , n3439 , n3441 );
or ( n3443 , n713 , n3311 , n3383 );
or ( n3444 , n3375 , n2796 );
nand ( n3445 , n3443 , n3444 );
nor ( n3446 , n3432 , n3442 , n3445 );
nand ( n3447 , n3363 , n3387 , n3423 , n3446 );
not ( n3448 , n3447 );
or ( n3449 , n2890 , n3448 );
and ( n3450 , n1317 , n2936 );
not ( n3451 , n1137 );
or ( n3452 , n2975 , n3451 );
not ( n3453 , n841 );
nand ( n3454 , n20 , n1408 );
not ( n3455 , n3454 );
or ( n3456 , n3453 , n3455 );
nand ( n3457 , n3456 , n1429 );
nand ( n3458 , n3452 , n3457 );
nor ( n3459 , n3450 , n3458 );
not ( n3460 , n1319 );
not ( n3461 , n3460 );
not ( n3462 , n2942 );
and ( n3463 , n3461 , n3462 );
and ( n3464 , n1730 , n2931 );
nor ( n3465 , n3463 , n3464 );
nand ( n3466 , n2996 , n1370 );
and ( n3467 , n1144 , n3012 );
and ( n3468 , n1419 , n2959 );
nor ( n3469 , n3467 , n3468 , n1403 );
and ( n3470 , n3008 , n1223 );
not ( n3471 , n1406 );
or ( n3472 , n3471 , n2950 );
not ( n3473 , n3015 );
or ( n3474 , n1612 , n3473 );
nand ( n3475 , n3472 , n3474 );
nor ( n3476 , n3470 , n3475 );
and ( n3477 , n3469 , n3476 );
nand ( n3478 , n3459 , n3465 , n3466 , n3477 );
and ( n3479 , n1852 , n3478 );
and ( n3480 , n1982 , n3108 );
nor ( n3481 , n3479 , n3480 );
nor ( n3482 , n2579 , n843 );
and ( n3483 , n3482 , n3033 );
and ( n3484 , n2018 , n3045 );
and ( n3485 , n2030 , n3059 );
nor ( n3486 , n3483 , n3484 , n3485 );
and ( n3487 , n2603 , n2916 );
not ( n3488 , n3064 );
and ( n3489 , n1985 , n3488 );
nor ( n3490 , n3487 , n3489 );
or ( n3491 , n841 , n2579 , n1411 );
and ( n3492 , n1998 , n3048 );
buf ( n3493 , n2781 );
not ( n3494 , n2324 );
nor ( n3495 , n3493 , n3494 );
not ( n3496 , n3495 );
nand ( n3497 , n1411 , n3496 );
and ( n3498 , n1849 , n3497 );
nor ( n3499 , n3492 , n3498 );
nand ( n3500 , n3491 , n3499 );
nand ( n3501 , n1982 , n2255 );
or ( n3502 , n3501 , n3041 );
not ( n3503 , n3078 );
or ( n3504 , n2015 , n3503 );
not ( n3505 , n16 );
not ( n3506 , n3505 );
not ( n3507 , n1992 );
and ( n3508 , n3506 , n3507 );
and ( n3509 , n1408 , n3069 );
nor ( n3510 , n3508 , n3509 );
or ( n3511 , n1411 , n3510 );
nand ( n3512 , n3502 , n3504 , n3511 );
nor ( n3513 , n3500 , n3512 );
and ( n3514 , n3481 , n3486 , n3490 , n3513 );
or ( n3515 , n2 , n3514 );
buf ( n3516 , n3493 );
or ( n3517 , n3516 , n3322 );
nand ( n3518 , n3517 , n713 );
and ( n3519 , n3384 , n3518 );
or ( n3520 , n2 , n11 );
not ( n3521 , n3520 );
or ( n3522 , n1980 , n3521 );
not ( n3523 , n1981 );
nand ( n3524 , n2 , n3523 );
nand ( n3525 , n3522 , n3524 );
and ( n3526 , n3525 , n3497 );
nor ( n3527 , n3519 , n3526 );
or ( n3528 , n3493 , n3134 );
nand ( n3529 , n3528 , n333 );
and ( n3530 , n80 , n3529 );
and ( n3531 , n2 , n1976 );
or ( n3532 , n3516 , n2330 );
nand ( n3533 , n3532 , n2412 );
and ( n3534 , n3531 , n3533 );
nor ( n3535 , n3530 , n3534 );
nand ( n3536 , n3515 , n3527 , n3535 );
nand ( n3537 , n3536 , n3 , n2299 );
nand ( n3538 , n3449 , n3537 );
and ( n3539 , n2526 , n3125 );
nor ( n3540 , n3539 , n841 , n2518 );
nor ( n3541 , n3538 , n3540 );
or ( n3542 , n2735 , n2378 );
and ( n3543 , n782 , n2371 );
nor ( n3544 , n3543 , n2473 );
or ( n3545 , n2518 , n3544 );
and ( n3546 , n2402 , n2679 , n2734 );
not ( n3547 , n2510 );
not ( n3548 , n20 );
nand ( n3549 , n3548 , n2517 );
nor ( n3550 , n3547 , n3549 );
not ( n3551 , n2851 );
and ( n3552 , n3550 , n3551 );
nor ( n3553 , n3546 , n3552 );
nand ( n3554 , n3542 , n3545 , n3553 );
not ( n3555 , n3550 );
not ( n3556 , n2540 );
not ( n3557 , n3556 );
or ( n3558 , n3555 , n3557 );
or ( n3559 , n2515 , n3278 );
nand ( n3560 , n3559 , n2734 , n2402 );
nand ( n3561 , n3558 , n3560 );
not ( n3562 , n2734 );
not ( n3563 , n3172 );
or ( n3564 , n3562 , n3563 );
nand ( n3565 , n415 , n3278 , n2519 );
nand ( n3566 , n3564 , n3565 );
nor ( n3567 , n3554 , n3561 , n3566 );
nand ( n3568 , n2572 , n2887 , n3541 , n3567 );
not ( n3569 , n4 );
nand ( n3570 , n3568 , n3569 );
nor ( n3571 , n963 , n2903 );
and ( n3572 , n3571 , n1424 );
not ( n3573 , n101 );
nor ( n3574 , n24 , n31 );
not ( n3575 , n3574 );
nand ( n3576 , n3573 , n3575 );
and ( n3577 , n3576 , n105 , n2900 );
nor ( n3578 , n910 , n3577 );
nor ( n3579 , n3572 , n3578 );
nor ( n3580 , n912 , n633 , n3577 );
not ( n3581 , n3580 );
and ( n3582 , n914 , n2922 );
nor ( n3583 , n910 , n2903 );
not ( n3584 , n3583 );
nor ( n3585 , n2084 , n3584 );
nor ( n3586 , n3582 , n3585 );
and ( n3587 , n3579 , n3581 , n3586 );
not ( n3588 , n3587 );
nor ( n3589 , n523 , n2903 );
and ( n3590 , n2512 , n3589 );
nor ( n3591 , n591 , n2903 );
and ( n3592 , n3591 , n2155 );
nor ( n3593 , n3590 , n3592 );
or ( n3594 , n2190 , n633 , n3577 );
nor ( n3595 , n571 , n2903 );
and ( n3596 , n3595 , n1882 );
nor ( n3597 , n585 , n3577 );
nor ( n3598 , n3596 , n3597 );
and ( n3599 , n3593 , n3594 , n3598 );
not ( n3600 , n3599 );
or ( n3601 , n3588 , n3600 );
nand ( n3602 , n3601 , n39 );
not ( n3603 , n17 );
not ( n3604 , n3575 );
and ( n3605 , n23 , n3604 );
not ( n3606 , n22 );
nor ( n3607 , n3605 , n3606 );
and ( n3608 , n39 , n3603 , n3607 );
not ( n3609 , n39 );
nor ( n3610 , n3609 , n692 );
not ( n3611 , n3610 );
nand ( n3612 , n3576 , n325 );
not ( n3613 , n3612 );
or ( n3614 , n3611 , n3613 );
or ( n3615 , n39 , n1411 );
nand ( n3616 , n3614 , n3615 );
nor ( n3617 , n3608 , n3616 );
not ( n3618 , n39 );
not ( n3619 , n2929 );
nor ( n3620 , n3619 , n910 );
or ( n3621 , n2924 , n913 );
not ( n3622 , n2959 );
or ( n3623 , n963 , n3622 );
nand ( n3624 , n3621 , n3623 );
nor ( n3625 , n3620 , n3624 );
not ( n3626 , n3625 );
and ( n3627 , n3618 , n3626 );
not ( n3628 , n20 );
nor ( n3629 , n3628 , n3609 );
and ( n3630 , n2935 , n3577 );
or ( n3631 , n2616 , n3630 );
or ( n3632 , n437 , n97 );
not ( n3633 , n3577 );
nand ( n3634 , n3632 , n3633 );
not ( n3635 , n2941 );
nand ( n3636 , n97 , n3635 );
and ( n3637 , n3634 , n2947 , n2949 , n3636 );
nand ( n3638 , n3631 , n3637 );
and ( n3639 , n3629 , n3638 );
nor ( n3640 , n3627 , n3639 );
and ( n3641 , n3602 , n3617 , n3640 );
not ( n3642 , n20 );
nor ( n3643 , n39 , n98 );
and ( n3644 , n3642 , n3643 , n2976 );
nand ( n3645 , n39 , n97 );
nor ( n3646 , n20 , n3645 );
not ( n3647 , n3646 );
nand ( n3648 , n3577 , n2974 );
not ( n3649 , n3648 );
or ( n3650 , n3647 , n3649 );
and ( n3651 , n1905 , n2615 , n2904 );
and ( n3652 , n2948 , n415 );
nor ( n3653 , n3651 , n3652 );
and ( n3654 , n2946 , n363 );
and ( n3655 , n438 , n2616 );
nor ( n3656 , n3655 , n3577 );
nor ( n3657 , n3654 , n3656 );
and ( n3658 , n3653 , n3657 );
nor ( n3659 , n3609 , n20 );
not ( n3660 , n3659 );
or ( n3661 , n3658 , n3660 );
nand ( n3662 , n3650 , n3661 );
nor ( n3663 , n3644 , n3662 );
nor ( n3664 , n39 , n2616 );
nand ( n3665 , n20 , n3664 , n2936 );
not ( n3666 , n20 );
not ( n3667 , n2952 );
or ( n3668 , n3666 , n3667 );
not ( n3669 , n3018 );
not ( n3670 , n20 );
and ( n3671 , n3669 , n3670 );
nor ( n3672 , n3671 , n39 );
nand ( n3673 , n3668 , n3672 );
nand ( n3674 , n584 , n2984 );
and ( n3675 , n1571 , n2993 );
and ( n3676 , n570 , n2987 );
nor ( n3677 , n3675 , n3676 );
and ( n3678 , n3674 , n3677 );
not ( n3679 , n3678 );
nand ( n3680 , n3679 , n3609 );
and ( n3681 , n3665 , n3673 , n3680 );
and ( n3682 , n3641 , n3663 , n3681 );
or ( n3683 , n3682 , n18 );
nand ( n3684 , n18 , n3609 );
or ( n3685 , n3684 , n3107 );
nor ( n3686 , n1984 , n98 );
nand ( n3687 , n3577 , n3058 );
nand ( n3688 , n39 , n3686 , n3687 );
nand ( n3689 , n3683 , n3685 , n3688 );
and ( n3690 , n584 , n2910 );
and ( n3691 , n766 , n2906 );
and ( n3692 , n782 , n2913 );
nor ( n3693 , n3690 , n3691 , n3692 );
or ( n3694 , n3684 , n3693 );
nand ( n3695 , n18 , n39 );
not ( n3696 , n2905 );
and ( n3697 , n766 , n3696 );
and ( n3698 , n3589 , n566 );
and ( n3699 , n3595 , n579 );
nor ( n3700 , n3698 , n3699 );
not ( n3701 , n3597 );
nand ( n3702 , n3700 , n3701 , n3594 );
nor ( n3703 , n3697 , n3702 );
or ( n3704 , n3695 , n3703 );
nor ( n3705 , n308 , n98 );
and ( n3706 , n3609 , n3705 , n3033 );
not ( n3707 , n3695 );
and ( n3708 , n3583 , n957 );
and ( n3709 , n3571 , n966 );
nor ( n3710 , n3708 , n3709 );
not ( n3711 , n3578 );
not ( n3712 , n3102 );
and ( n3713 , n914 , n3712 );
nor ( n3714 , n3713 , n3580 );
nand ( n3715 , n3710 , n3711 , n3714 );
and ( n3716 , n3707 , n3715 );
nor ( n3717 , n3706 , n3716 );
nand ( n3718 , n3694 , n3704 , n3717 );
or ( n3719 , n2862 , n1316 , n39 , n3503 );
nand ( n3720 , n3577 , n3040 );
and ( n3721 , n2615 , n3720 );
and ( n3722 , n2948 , n859 );
and ( n3723 , n2946 , n366 );
nor ( n3724 , n434 , n3577 );
nor ( n3725 , n3722 , n3723 , n3724 );
not ( n3726 , n3725 );
nor ( n3727 , n3721 , n3726 );
or ( n3728 , n3660 , n3727 );
nand ( n3729 , n3728 , n3617 );
nand ( n3730 , n18 , n3729 );
and ( n3731 , n3609 , n1582 , n3065 );
nand ( n3732 , n3577 , n3032 );
and ( n3733 , n39 , n3705 , n3732 );
nor ( n3734 , n3731 , n3733 );
nor ( n3735 , n20 , n39 );
and ( n3736 , n18 , n3735 , n3052 );
and ( n3737 , n3577 , n3077 );
or ( n3738 , n2616 , n3737 );
not ( n3739 , n3063 );
not ( n3740 , n3062 );
nor ( n3741 , n3739 , n3724 , n3740 );
nand ( n3742 , n3738 , n3741 );
and ( n3743 , n39 , n1582 , n3742 );
nor ( n3744 , n3736 , n3743 );
nand ( n3745 , n3719 , n3730 , n3734 , n3744 );
nor ( n3746 , n3689 , n3718 , n3745 );
or ( n3747 , n1848 , n3520 );
buf ( n3748 , n3747 );
or ( n3749 , n2299 , n4 );
nor ( n3750 , n3 , n3749 );
nand ( n3751 , n1 , n3750 );
nor ( n3752 , n3746 , n3748 , n3751 );
and ( n3753 , n4 , n2299 );
and ( n3754 , n2298 , n3753 );
nand ( n3755 , n1 , n3754 );
nor ( n3756 , n11 , n13 );
or ( n3757 , n12 , n3756 );
not ( n3758 , n2 );
nand ( n3759 , n3757 , n3758 );
and ( n3760 , n38 , n3609 );
not ( n3761 , n3760 );
not ( n3762 , n3761 );
not ( n3763 , n3762 );
not ( n3764 , n3763 );
not ( n3765 , n3764 );
not ( n3766 , n3765 );
not ( n3767 , n3766 );
not ( n3768 , n3767 );
not ( n3769 , n3768 );
and ( n3770 , n3769 , n3495 );
nor ( n3771 , n3493 , n3765 );
nand ( n3772 , n3576 , n2327 );
and ( n3773 , n3771 , n3772 );
not ( n3774 , n17 );
and ( n3775 , n92 , n3764 , n3612 );
and ( n3776 , n3765 , n703 );
nor ( n3777 , n3775 , n3776 );
or ( n3778 , n3774 , n3777 );
or ( n3779 , n22 , n3764 );
or ( n3780 , n3763 , n3607 );
not ( n3781 , n17 );
nand ( n3782 , n3779 , n3780 , n3781 );
nand ( n3783 , n3778 , n3782 );
nor ( n3784 , n3770 , n3773 , n3783 );
or ( n3785 , n3759 , n3784 );
not ( n3786 , n3747 );
and ( n3787 , n18 , n3786 );
nand ( n3788 , n454 , n3787 );
not ( n3789 , n2349 );
not ( n3790 , n3789 );
not ( n3791 , n3777 );
and ( n3792 , n3790 , n3791 );
nor ( n3793 , n14 , n3782 );
nor ( n3794 , n3792 , n3793 );
or ( n3795 , n3788 , n3794 );
not ( n3796 , n78 );
not ( n3797 , n3796 );
nor ( n3798 , n38 , n3797 );
not ( n3799 , n13 );
and ( n3800 , n1980 , n3799 );
and ( n3801 , n3800 , n3529 );
not ( n3802 , n1848 );
not ( n3803 , n3802 );
not ( n3804 , n3803 );
and ( n3805 , n3804 , n3334 );
nor ( n3806 , n3801 , n3805 );
not ( n3807 , n3806 );
and ( n3808 , n3798 , n3807 );
not ( n3809 , n3803 );
not ( n3810 , n3809 );
and ( n3811 , n17 , n3493 );
nand ( n3812 , n23 , n31 );
not ( n3813 , n3812 );
nand ( n3814 , n22 , n3813 );
not ( n3815 , n3814 );
and ( n3816 , n40 , n3815 );
not ( n3817 , n40 );
not ( n3818 , n22 );
nand ( n3819 , n23 , n24 );
or ( n3820 , n31 , n3819 );
or ( n3821 , n3818 , n3820 );
nand ( n3822 , n3814 , n3821 );
and ( n3823 , n3817 , n3822 );
nor ( n3824 , n3816 , n3823 );
nor ( n3825 , n3811 , n3824 );
not ( n3826 , n17 );
not ( n3827 , n563 );
nand ( n3828 , n3826 , n3827 );
not ( n3829 , n3828 );
nor ( n3830 , n3493 , n2327 );
nor ( n3831 , n3825 , n3829 , n3830 );
nand ( n3832 , n38 , n3796 );
nor ( n3833 , n3810 , n39 , n3831 , n3832 );
nor ( n3834 , n3808 , n3833 );
nand ( n3835 , n3785 , n3795 , n3834 );
not ( n3836 , n38 );
nand ( n3837 , n12 , n13 );
nand ( n3838 , n3837 , n1981 );
not ( n3839 , n3838 );
nand ( n3840 , n2 , n3836 , n3839 , n3533 );
not ( n3841 , n20 );
nand ( n3842 , n3841 , n3767 );
not ( n3843 , n3842 );
nand ( n3844 , n3843 , n3787 );
not ( n3845 , n3844 );
nand ( n3846 , n3845 , n3033 , n97 );
nor ( n3847 , n308 , n3748 );
nand ( n3848 , n38 , n3847 , n3643 , n3732 );
not ( n3849 , n455 );
nand ( n3850 , n3766 , n3849 );
not ( n3851 , n3850 );
nand ( n3852 , n3851 , n3787 , n3720 );
nand ( n3853 , n3840 , n3846 , n3848 , n3852 );
not ( n3854 , n2 );
or ( n3855 , n3854 , n3839 , n3784 );
and ( n3856 , n39 , n2341 );
nor ( n3857 , n445 , n39 );
not ( n3858 , n3857 );
not ( n3859 , n17 );
not ( n3860 , n40 );
nand ( n3861 , n3860 , n3815 );
nand ( n3862 , n40 , n3822 );
nand ( n3863 , n3861 , n276 , n3862 );
and ( n3864 , n3859 , n3863 );
not ( n3865 , n3863 );
not ( n3866 , n2323 );
and ( n3867 , n3865 , n3866 );
nor ( n3868 , n3867 , n1891 );
and ( n3869 , n325 , n3861 , n3862 );
nor ( n3870 , n3869 , n692 );
nor ( n3871 , n3864 , n3868 , n3870 );
or ( n3872 , n3858 , n3871 );
not ( n3873 , n2781 );
nand ( n3874 , n39 , n3873 );
or ( n3875 , n3874 , n2330 );
nand ( n3876 , n3872 , n3875 );
not ( n3877 , n3610 );
nor ( n3878 , n3877 , n2353 );
nor ( n3879 , n3856 , n3876 , n3878 );
nor ( n3880 , n39 , n2781 );
nand ( n3881 , n445 , n3880 , n3772 );
nor ( n3882 , n17 , n39 );
nand ( n3883 , n445 , n3882 , n3607 );
nand ( n3884 , n3609 , n445 , n693 , n3612 );
nand ( n3885 , n3879 , n3881 , n3883 , n3884 );
nand ( n3886 , n2 , n38 , n3839 , n3885 );
nand ( n3887 , n3855 , n3886 );
nand ( n3888 , n325 , n3824 );
nand ( n3889 , n3802 , n693 , n3609 , n3888 );
not ( n3890 , n3889 );
not ( n3891 , n17 );
nand ( n3892 , n3857 , n3800 , n3891 , n3607 );
and ( n3893 , n2112 , n39 , n3800 );
and ( n3894 , n39 , n3802 , n711 );
nor ( n3895 , n3893 , n3894 );
not ( n3896 , n3516 );
nand ( n3897 , n3896 , n3800 , n3857 , n3772 );
not ( n3898 , n3874 );
and ( n3899 , n3266 , n3800 , n3898 );
not ( n3900 , n3800 );
nor ( n3901 , n3900 , n39 , n41 , n3871 );
nor ( n3902 , n3899 , n3901 );
nand ( n3903 , n3892 , n3895 , n3897 , n3902 );
nand ( n3904 , n39 , n3800 );
or ( n3905 , n3904 , n319 );
nand ( n3906 , n3857 , n3800 , n693 , n3612 );
not ( n3907 , n40 );
nor ( n3908 , n3609 , n3907 );
nand ( n3909 , n3908 , n693 , n3802 , n326 );
nand ( n3910 , n3905 , n3906 , n3909 );
not ( n3911 , n3610 );
not ( n3912 , n702 );
not ( n3913 , n40 );
nand ( n3914 , n3913 , n13 );
nor ( n3915 , n3911 , n12 , n3912 , n3914 );
nor ( n3916 , n3890 , n3903 , n3910 , n3915 );
or ( n3917 , n3832 , n3916 );
not ( n3918 , n3322 );
not ( n3919 , n3769 );
not ( n3920 , n3919 );
nor ( n3921 , n3516 , n3797 );
nand ( n3922 , n3918 , n3920 , n3809 , n3921 );
nand ( n3923 , n3917 , n3922 );
or ( n3924 , n3835 , n3853 , n3887 , n3923 );
or ( n3925 , n3844 , n3051 );
and ( n3926 , n3783 , n2733 , n3787 );
nand ( n3927 , n38 , n3735 );
not ( n3928 , n3787 );
nor ( n3929 , n3725 , n3927 , n3928 );
nor ( n3930 , n3926 , n3929 );
nand ( n3931 , n3847 , n306 , n3783 );
nand ( n3932 , n3925 , n3930 , n3931 );
not ( n3933 , n3693 );
not ( n3934 , n3766 );
not ( n3935 , n3934 );
not ( n3936 , n3935 );
not ( n3937 , n3936 );
not ( n3938 , n3937 );
and ( n3939 , n3933 , n3938 , n3787 );
and ( n3940 , n3591 , n621 );
nor ( n3941 , n3940 , n3702 );
or ( n3942 , n3928 , n3938 , n3941 );
nor ( n3943 , n3766 , n455 );
not ( n3944 , n3943 );
or ( n3945 , n3041 , n3928 , n3944 );
nand ( n3946 , n3942 , n3945 );
nor ( n3947 , n3939 , n3946 );
not ( n3948 , n2067 );
not ( n3949 , n3794 );
and ( n3950 , n3948 , n3949 );
and ( n3951 , n2110 , n3783 );
nor ( n3952 , n3950 , n3951 );
and ( n3953 , n3920 , n3106 );
not ( n3954 , n3936 );
and ( n3955 , n3954 , n3715 );
nor ( n3956 , n3953 , n3955 );
nand ( n3957 , n3952 , n3956 );
nand ( n3958 , n20 , n3766 );
or ( n3959 , n3958 , n3741 );
nand ( n3960 , n3935 , n2068 );
not ( n3961 , n3960 );
not ( n3962 , n3737 );
and ( n3963 , n3961 , n3962 );
not ( n3964 , n2068 );
nor ( n3965 , n3935 , n3964 );
and ( n3966 , n3965 , n3078 );
nor ( n3967 , n3963 , n3966 );
nor ( n3968 , n3767 , n98 );
and ( n3969 , n20 , n3968 , n3687 );
not ( n3970 , n20 );
nor ( n3971 , n3970 , n3768 );
and ( n3972 , n3971 , n3065 );
nor ( n3973 , n3969 , n3972 );
nand ( n3974 , n3959 , n3967 , n3973 );
or ( n3975 , n3957 , n3974 );
nand ( n3976 , n3975 , n3787 );
or ( n3977 , n3937 , n3625 );
not ( n3978 , n3958 );
not ( n3979 , n3637 );
and ( n3980 , n3978 , n3979 );
and ( n3981 , n3965 , n2936 );
nor ( n3982 , n3980 , n3981 );
nand ( n3983 , n3977 , n3982 , n3952 );
or ( n3984 , n3920 , n3587 );
not ( n3985 , n3971 );
or ( n3986 , n3985 , n2952 );
or ( n3987 , n3960 , n3630 );
nand ( n3988 , n3984 , n3986 , n3987 );
or ( n3989 , n3983 , n3988 );
nor ( n3990 , n18 , n3747 );
nand ( n3991 , n3989 , n3990 );
not ( n3992 , n3937 );
or ( n3993 , n3992 , n3599 );
or ( n3994 , n3927 , n3658 );
and ( n3995 , n3648 , n3935 , n2573 );
and ( n3996 , n3843 , n3018 );
nor ( n3997 , n3995 , n3996 );
nand ( n3998 , n3993 , n3994 , n3997 );
not ( n3999 , n2237 );
not ( n4000 , n3783 );
or ( n4001 , n3999 , n4000 );
nand ( n4002 , n2976 , n3920 , n2573 );
nand ( n4003 , n4001 , n4002 );
or ( n4004 , n3678 , n3954 );
or ( n4005 , n2261 , n3777 );
or ( n4006 , n2242 , n3782 );
nand ( n4007 , n4004 , n4005 , n4006 );
or ( n4008 , n3998 , n4003 , n4007 );
nand ( n4009 , n4008 , n3990 );
nand ( n4010 , n3947 , n3976 , n3991 , n4009 );
nor ( n4011 , n3924 , n3932 , n4010 );
or ( n4012 , n3755 , n4011 );
and ( n4013 , n3836 , n3609 );
not ( n4014 , n4013 );
not ( n4015 , n4014 );
not ( n4016 , n4015 );
not ( n4017 , n4016 );
not ( n4018 , n4017 );
not ( n4019 , n4018 );
nor ( n4020 , n20 , n4019 );
and ( n4021 , n3052 , n4020 , n3787 );
not ( n4022 , n14 );
or ( n4023 , n22 , n4017 );
or ( n4024 , n4016 , n3607 );
not ( n4025 , n17 );
nand ( n4026 , n4023 , n4024 , n4025 );
not ( n4027 , n4026 );
not ( n4028 , n4027 );
or ( n4029 , n4022 , n4028 );
and ( n4030 , n92 , n4017 , n3612 );
and ( n4031 , n4018 , n703 );
nor ( n4032 , n4030 , n4031 );
or ( n4033 , n2244 , n4032 );
nand ( n4034 , n4029 , n4033 );
and ( n4035 , n2066 , n4034 );
not ( n4036 , n2649 );
not ( n4037 , n17 );
or ( n4038 , n4037 , n4032 );
nand ( n4039 , n4038 , n4026 );
not ( n4040 , n4039 );
or ( n4041 , n4036 , n4040 );
nand ( n4042 , n908 , n4039 );
nand ( n4043 , n4041 , n4042 );
nor ( n4044 , n4035 , n4043 );
not ( n4045 , n4019 );
not ( n4046 , n4045 );
not ( n4047 , n4046 );
not ( n4048 , n4047 );
not ( n4049 , n4048 );
and ( n4050 , n4049 , n3106 );
not ( n4051 , n4049 );
and ( n4052 , n4051 , n3715 );
nor ( n4053 , n4050 , n4052 );
nor ( n4054 , n4045 , n2629 );
and ( n4055 , n4054 , n3687 );
nor ( n4056 , n4046 , n2629 );
and ( n4057 , n4056 , n3059 );
nor ( n4058 , n4055 , n4057 );
nand ( n4059 , n20 , n4019 );
not ( n4060 , n4059 );
and ( n4061 , n4060 , n3742 );
not ( n4062 , n20 );
nor ( n4063 , n4062 , n4048 );
or ( n4064 , n2616 , n3503 );
nand ( n4065 , n4064 , n3064 );
and ( n4066 , n4063 , n4065 );
nor ( n4067 , n4061 , n4066 );
nand ( n4068 , n4044 , n4053 , n4058 , n4067 );
and ( n4069 , n3787 , n4068 );
nor ( n4070 , n4021 , n4069 );
not ( n4071 , n4070 );
nand ( n4072 , n3809 , n3798 );
or ( n4073 , n4072 , n39 , n3831 );
not ( n4074 , n2600 );
nand ( n4075 , n3847 , n4074 , n4039 );
nand ( n4076 , n4073 , n4075 );
or ( n4077 , n3832 , n3806 );
not ( n4078 , n3788 );
nand ( n4079 , n4078 , n4034 );
nand ( n4080 , n4077 , n4079 );
not ( n4081 , n4049 );
buf ( n4082 , n4081 );
not ( n4083 , n4082 );
or ( n4084 , n3703 , n4083 , n3928 );
nor ( n4085 , n4019 , n2230 );
nand ( n4086 , n3033 , n3787 , n4085 );
nand ( n4087 , n4084 , n4086 );
nor ( n4088 , n4071 , n4076 , n4080 , n4087 );
not ( n4089 , n3916 );
and ( n4090 , n3798 , n4089 );
nand ( n4091 , n3836 , n3735 );
or ( n4092 , n3727 , n4091 , n3928 );
nor ( n4093 , n4045 , n2230 );
nand ( n4094 , n4093 , n3787 , n3732 );
nand ( n4095 , n4092 , n4094 );
not ( n4096 , n4083 );
nor ( n4097 , n3693 , n4096 , n3928 );
nor ( n4098 , n4090 , n4095 , n4097 );
not ( n4099 , n3759 );
not ( n4100 , n4081 );
and ( n4101 , n4100 , n3495 );
and ( n4102 , n3836 , n3880 );
and ( n4103 , n4102 , n3772 );
nor ( n4104 , n4101 , n4103 , n4039 );
not ( n4105 , n4104 );
and ( n4106 , n4099 , n4105 );
nand ( n4107 , n2195 , n4039 );
nor ( n4108 , n3928 , n4107 );
nor ( n4109 , n4106 , n4108 );
not ( n4110 , n3322 );
nand ( n4111 , n4110 , n3809 , n4083 , n3921 );
nand ( n4112 , n4039 , n305 , n2440 );
nor ( n4113 , n3630 , n4059 );
nand ( n4114 , n4113 , n2816 , n450 );
and ( n4115 , n4112 , n4042 , n4114 );
not ( n4116 , n4032 );
not ( n4117 , n3789 );
nand ( n4118 , n4116 , n4117 , n2066 );
not ( n4119 , n3625 );
and ( n4120 , n4119 , n4100 );
and ( n4121 , n2549 , n4027 );
nor ( n4122 , n4120 , n4121 );
nand ( n4123 , n4115 , n4118 , n4122 );
not ( n4124 , n4063 );
and ( n4125 , n2936 , n2816 , n450 );
nor ( n4126 , n4125 , n2951 );
or ( n4127 , n4124 , n4126 );
or ( n4128 , n3587 , n4100 );
or ( n4129 , n4059 , n3637 );
nand ( n4130 , n4127 , n4128 , n4129 );
or ( n4131 , n4123 , n4130 );
nand ( n4132 , n4131 , n3990 );
or ( n4133 , n4081 , n3678 );
nor ( n4134 , n20 , n2600 );
nand ( n4135 , n4134 , n4039 );
and ( n4136 , n4093 , n3648 );
and ( n4137 , n454 , n4034 );
nor ( n4138 , n4136 , n4137 );
nand ( n4139 , n4133 , n4135 , n4107 , n4138 );
not ( n4140 , n4082 );
or ( n4141 , n4140 , n3599 );
or ( n4142 , n3658 , n4091 );
and ( n4143 , n4020 , n3018 );
and ( n4144 , n4085 , n2976 );
nor ( n4145 , n4143 , n4144 );
nand ( n4146 , n4141 , n4142 , n4145 );
or ( n4147 , n4139 , n4146 );
nand ( n4148 , n4147 , n3990 );
and ( n4149 , n4111 , n4132 , n4148 );
and ( n4150 , n4088 , n4098 , n4109 , n4149 );
nand ( n4151 , n2506 , n3750 );
or ( n4152 , n4150 , n4151 );
nand ( n4153 , n4012 , n4152 );
nor ( n4154 , n3752 , n4153 );
nor ( n4155 , n41 , n3749 , n3838 );
nand ( n4156 , n1 , n2298 );
not ( n4157 , n4156 );
and ( n4158 , n2 , n4157 );
not ( n4159 , n4158 );
nor ( n4160 , n3609 , n4159 );
not ( n4161 , n325 );
and ( n4162 , n693 , n4161 );
nor ( n4163 , n4162 , n3830 );
nand ( n4164 , n4163 , n3828 , n3576 );
and ( n4165 , n4155 , n4160 , n4164 );
not ( n4166 , n3749 );
nand ( n4167 , n3609 , n4166 );
or ( n4168 , n4159 , n4167 , n3838 );
nand ( n4169 , n38 , n2508 );
or ( n4170 , n4169 , n3749 , n1971 );
nand ( n4171 , n4168 , n4170 );
and ( n4172 , n4171 , n3533 );
nor ( n4173 , n4165 , n4172 );
nand ( n4174 , n5 , n3836 );
nor ( n4175 , n4 , n4174 , n1971 );
and ( n4176 , n4175 , n2508 , n3885 );
not ( n4177 , n3384 );
nor ( n4178 , n4177 , n3751 );
and ( n4179 , n3609 , n4178 , n3518 );
nor ( n4180 , n4176 , n4179 );
and ( n4181 , n4173 , n4180 );
and ( n4182 , n1 , n3 );
not ( n4183 , n4182 );
nor ( n4184 , n2506 , n5 );
nand ( n4185 , n4183 , n4184 );
or ( n4186 , n3569 , n4185 );
nor ( n4187 , n2298 , n2299 );
or ( n4188 , n4 , n4187 );
nand ( n4189 , n4186 , n4188 , n3536 );
nand ( n4190 , n3570 , n4154 , n4181 , n4189 );
and ( n4191 , n1845 , n3800 );
not ( n4192 , n1851 );
nor ( n4193 , n4191 , n4192 );
nor ( n4194 , n4193 , n3749 , n4159 );
or ( n4195 , n39 , n3496 );
not ( n4196 , n3772 );
or ( n4197 , n3874 , n4196 );
nand ( n4198 , n4195 , n4197 , n3617 );
and ( n4199 , n4194 , n4198 );
nand ( n4200 , n4166 , n2508 );
or ( n4201 , n4200 , n4193 , n4104 );
not ( n4202 , n4198 );
or ( n4203 , n4202 , n3759 , n3751 );
nand ( n4204 , n4201 , n4203 );
not ( n4205 , n13 );
nor ( n4206 , n3118 , n3751 );
nand ( n4207 , n39 , n445 , n4205 , n4206 );
nor ( n4208 , n3609 , n445 );
nand ( n4209 , n4208 , n4158 , n4166 , n3839 );
and ( n4210 , n4207 , n4209 );
nor ( n4211 , n4210 , n3871 );
nor ( n4212 , n4199 , n4204 , n4211 );
and ( n4213 , n3888 , n3610 , n4178 );
nand ( n4214 , n39 , n3370 );
nor ( n4215 , n3831 , n3751 , n4214 );
nor ( n4216 , n4213 , n4215 );
not ( n4217 , n13 );
nand ( n4218 , n4208 , n4206 , n4217 , n4164 );
not ( n4219 , n13 );
nand ( n4220 , n4219 , n3609 , n4206 , n3529 );
nand ( n4221 , n4212 , n4216 , n4218 , n4220 );
or ( n4222 , n4190 , n4221 );
nor ( n4223 , n6 , n7 );
not ( n4224 , n4223 );
not ( n4225 , n4224 );
buf ( n4226 , n4225 );
not ( n4227 , n4226 );
not ( n4228 , n4227 );
not ( n4229 , n4228 );
not ( n4230 , n4229 );
not ( n4231 , n4230 );
not ( n4232 , n4231 );
not ( n4233 , n4232 );
not ( n4234 , n9 );
not ( n4235 , n8 );
not ( n4236 , n10 );
and ( n4237 , n4234 , n4235 , n4236 );
nor ( n4238 , n4233 , n4237 );
nand ( n4239 , n4222 , n4238 );
nand ( n4240 , n3569 , n2300 );
not ( n4241 , n4240 );
and ( n4242 , n4223 , n4237 );
not ( n4243 , n4242 );
nor ( n4244 , n2 , n4241 , n4243 );
not ( n4245 , n3514 );
and ( n4246 , n4244 , n4245 );
not ( n4247 , n2051 );
not ( n4248 , n2 );
and ( n4249 , n1 , n4223 );
nor ( n4250 , n4 , n5 );
not ( n4251 , n4250 );
not ( n4252 , n4251 );
not ( n4253 , n4252 );
nor ( n4254 , n3 , n4253 );
nand ( n4255 , n4248 , n4237 , n4249 , n4254 );
nor ( n4256 , n4247 , n4255 );
nor ( n4257 , n4246 , n4256 );
nor ( n4258 , n4231 , n4241 );
and ( n4259 , n4258 , n3520 , n4237 );
and ( n4260 , n4259 , n3497 );
not ( n4261 , n4232 );
not ( n4262 , n4261 );
not ( n4263 , n4262 );
and ( n4264 , n22 , n4263 );
not ( n4265 , n4251 );
and ( n4266 , n4265 , n4242 );
nand ( n4267 , n4266 , n3520 , n2507 );
not ( n4268 , n2884 );
or ( n4269 , n4267 , n4268 );
not ( n4270 , n4266 );
nor ( n4271 , n4270 , n4156 , n3521 );
not ( n4272 , n1842 );
nand ( n4273 , n4271 , n4272 );
nand ( n4274 , n4269 , n4273 );
nor ( n4275 , n4260 , n4264 , n4274 );
not ( n4276 , n2 );
and ( n4277 , n2506 , n4276 , n4254 , n4242 );
nand ( n4278 , n4277 , n3113 );
nand ( n4279 , n4239 , n4257 , n4275 , n4278 );
not ( n4280 , n4255 );
not ( n4281 , n18 );
and ( n4282 , n23 , n4281 , n3256 );
not ( n4283 , n23 );
nor ( n4284 , n4283 , n1409 );
nor ( n4285 , n4282 , n4284 );
not ( n4286 , n348 );
nor ( n4287 , n27 , n28 );
buf ( n4288 , n4287 );
or ( n4289 , n25 , n4288 );
and ( n4290 , n4286 , n4289 );
nand ( n4291 , n32 , n4290 );
buf ( n4292 , n4291 );
not ( n4293 , n4292 );
not ( n4294 , n25 );
not ( n4295 , n27 );
nand ( n4296 , n4295 , n30 );
nor ( n4297 , n27 , n28 );
nand ( n4298 , n4296 , n4297 );
buf ( n4299 , n4298 );
buf ( n4300 , n4299 );
not ( n4301 , n4300 );
not ( n4302 , n4301 );
not ( n4303 , n4302 );
or ( n4304 , n4294 , n4303 );
not ( n4305 , n4288 );
not ( n4306 , n4305 );
not ( n4307 , n4306 );
and ( n4308 , n234 , n4307 );
not ( n4309 , n22 );
not ( n4310 , n23 );
nand ( n4311 , n4309 , n4310 );
nand ( n4312 , n998 , n4311 );
nand ( n4313 , n998 , n4312 );
not ( n4314 , n4313 );
buf ( n4315 , n4314 );
not ( n4316 , n4315 );
nor ( n4317 , n4308 , n4316 );
nand ( n4318 , n4304 , n4317 );
not ( n4319 , n4318 );
not ( n4320 , n4319 );
or ( n4321 , n4293 , n4320 );
not ( n4322 , n4316 );
buf ( n4323 , n4322 );
not ( n4324 , n4302 );
nand ( n4325 , n4323 , n1382 , n4324 );
nand ( n4326 , n4321 , n4325 );
and ( n4327 , n1419 , n4326 );
not ( n4328 , n16 );
not ( n4329 , n23 );
nor ( n4330 , n4328 , n4329 );
and ( n4331 , n4330 , n1958 );
nor ( n4332 , n4327 , n4331 );
not ( n4333 , n26 );
nor ( n4334 , n4333 , n32 );
nor ( n4335 , n25 , n4288 );
not ( n4336 , n4335 );
not ( n4337 , n4336 );
nand ( n4338 , n4334 , n4337 );
not ( n4339 , n32 );
not ( n4340 , n26 );
not ( n4341 , n4340 );
nor ( n4342 , n25 , n37 );
not ( n4343 , n4342 );
or ( n4344 , n4341 , n4343 );
not ( n4345 , n32 );
nand ( n4346 , n4344 , n4345 );
not ( n4347 , n4346 );
or ( n4348 , n4339 , n4347 );
not ( n4349 , n26 );
not ( n4350 , n26 );
nand ( n4351 , n4350 , n25 );
nand ( n4352 , n4349 , n4351 );
not ( n4353 , n4287 );
nand ( n4354 , n232 , n4353 );
nor ( n4355 , n4352 , n4354 );
nand ( n4356 , n4348 , n4355 );
not ( n4357 , n4356 );
not ( n4358 , n4357 );
and ( n4359 , n4338 , n4358 );
not ( n4360 , n4300 );
not ( n4361 , n166 );
not ( n4362 , n177 );
nand ( n4363 , n391 , n4361 , n4362 );
nand ( n4364 , n4360 , n4363 );
not ( n4365 , n4364 );
not ( n4366 , n4365 );
nand ( n4367 , n25 , n26 );
nor ( n4368 , n32 , n4367 );
not ( n4369 , n4368 );
not ( n4370 , n26 );
not ( n4371 , n4288 );
nor ( n4372 , n32 , n37 );
nand ( n4373 , n4371 , n4372 );
nand ( n4374 , n4373 , n4346 );
nand ( n4375 , n4370 , n4374 );
nand ( n4376 , n4369 , n4375 );
nand ( n4377 , n4366 , n4376 );
nand ( n4378 , n4359 , n4377 );
not ( n4379 , n4313 );
not ( n4380 , n4379 );
nor ( n4381 , n4337 , n4380 );
not ( n4382 , n4381 );
not ( n4383 , n4365 );
or ( n4384 , n4382 , n4383 );
buf ( n4385 , n27 );
or ( n4386 , n28 , n25 , n4385 );
nand ( n4387 , n4386 , n32 );
nand ( n4388 , n4387 , n4379 );
buf ( n4389 , n4388 );
nand ( n4390 , n4384 , n4389 );
and ( n4391 , n4292 , n4390 );
not ( n4392 , n22 );
and ( n4393 , n4392 , n1094 );
not ( n4394 , n4366 );
and ( n4395 , n4393 , n4394 );
nor ( n4396 , n4391 , n4395 );
or ( n4397 , n4378 , n4396 );
not ( n4398 , n4397 );
and ( n4399 , n1940 , n4398 );
and ( n4400 , n4330 , n1314 );
nor ( n4401 , n4399 , n4400 );
not ( n4402 , n4359 );
not ( n4403 , n4376 );
not ( n4404 , n389 );
not ( n4405 , n4299 );
nand ( n4406 , n4404 , n4405 );
and ( n4407 , n34 , n4406 );
not ( n4408 , n34 );
not ( n4409 , n4408 );
not ( n4410 , n4299 );
or ( n4411 , n4409 , n4410 );
nand ( n4412 , n4411 , n4363 );
nor ( n4413 , n4407 , n4412 );
buf ( n4414 , n4413 );
nor ( n4415 , n4403 , n4414 );
nor ( n4416 , n4402 , n4415 );
not ( n4417 , n4416 );
not ( n4418 , n4315 );
nor ( n4419 , n4337 , n4418 );
not ( n4420 , n4419 );
not ( n4421 , n4414 );
or ( n4422 , n4420 , n4421 );
nand ( n4423 , n4422 , n4389 );
and ( n4424 , n4292 , n4423 );
and ( n4425 , n4393 , n4414 );
nor ( n4426 , n4424 , n4425 );
nor ( n4427 , n4417 , n4426 );
not ( n4428 , n4427 );
not ( n4429 , n4428 );
and ( n4430 , n1613 , n4429 );
not ( n4431 , n1947 );
not ( n4432 , n32 );
not ( n4433 , n26 );
not ( n4434 , n4433 );
not ( n4435 , n475 );
or ( n4436 , n4434 , n4435 );
not ( n4437 , n32 );
nand ( n4438 , n4436 , n4437 );
not ( n4439 , n4438 );
or ( n4440 , n4432 , n4439 );
nand ( n4441 , n37 , n4353 );
nor ( n4442 , n4352 , n4441 );
nand ( n4443 , n4440 , n4442 );
buf ( n4444 , n4443 );
not ( n4445 , n4444 );
not ( n4446 , n4445 );
nand ( n4447 , n4338 , n4446 );
not ( n4448 , n26 );
not ( n4449 , n605 );
not ( n4450 , n4449 );
not ( n4451 , n4305 );
or ( n4452 , n4450 , n4451 );
nand ( n4453 , n4452 , n4438 );
nand ( n4454 , n4448 , n4453 );
not ( n4455 , n4454 );
nor ( n4456 , n4368 , n4455 );
and ( n4457 , n391 , n190 , n384 );
not ( n4458 , n4457 );
nor ( n4459 , n4385 , n28 );
nand ( n4460 , n4458 , n4459 , n4296 );
not ( n4461 , n4460 );
nor ( n4462 , n4456 , n4461 );
nor ( n4463 , n4447 , n4462 );
not ( n4464 , n4291 );
buf ( n4465 , n4289 );
nand ( n4466 , n4465 , n4379 );
not ( n4467 , n4299 );
nor ( n4468 , n34 , n36 );
and ( n4469 , n190 , n4468 );
nand ( n4470 , n391 , n4469 );
nand ( n4471 , n4467 , n4470 );
or ( n4472 , n4466 , n4471 );
nand ( n4473 , n4472 , n4388 );
not ( n4474 , n4473 );
or ( n4475 , n4464 , n4474 );
not ( n4476 , n4393 );
or ( n4477 , n4476 , n4471 );
nand ( n4478 , n4475 , n4477 );
nand ( n4479 , n4463 , n4478 );
not ( n4480 , n4479 );
and ( n4481 , n4431 , n4480 );
nor ( n4482 , n4430 , n4481 );
and ( n4483 , n4285 , n4332 , n4401 , n4482 );
or ( n4484 , n22 , n1021 );
not ( n4485 , n4484 );
not ( n4486 , n32 );
and ( n4487 , n4486 , n4314 );
nand ( n4488 , n35 , n4487 );
not ( n4489 , n4488 );
not ( n4490 , n160 );
not ( n4491 , n29 );
nand ( n4492 , n4491 , n34 );
not ( n4493 , n4298 );
nand ( n4494 , n4492 , n4493 );
nor ( n4495 , n4457 , n4494 );
not ( n4496 , n4495 );
not ( n4497 , n4496 );
not ( n4498 , n4497 );
not ( n4499 , n4498 );
or ( n4500 , n4490 , n4499 );
not ( n4501 , n4494 );
not ( n4502 , n4501 );
and ( n4503 , n199 , n4502 );
nor ( n4504 , n4503 , n4337 );
nand ( n4505 , n4500 , n4504 );
not ( n4506 , n4505 );
nand ( n4507 , n4323 , n4506 );
not ( n4508 , n4507 );
or ( n4509 , n4489 , n4508 );
not ( n4510 , n26 );
not ( n4511 , n4471 );
buf ( n4512 , n4492 );
nand ( n4513 , n4511 , n4512 );
not ( n4514 , n4513 );
nand ( n4515 , n1053 , n4453 );
buf ( n4516 , n4443 );
and ( n4517 , n4515 , n4516 );
nand ( n4518 , n4510 , n4514 , n4517 );
not ( n4519 , n4515 );
not ( n4520 , n4519 );
not ( n4521 , n4445 );
nand ( n4522 , n4506 , n4520 , n4514 , n4521 );
not ( n4523 , n2315 );
not ( n4524 , n1075 );
nand ( n4525 , n4523 , n4524 );
not ( n4526 , n4525 );
not ( n4527 , n4526 );
not ( n4528 , n4527 );
not ( n4529 , n4497 );
and ( n4530 , n4528 , n4529 );
not ( n4531 , n1000 );
nand ( n4532 , n4531 , n4335 );
not ( n4533 , n4532 );
not ( n4534 , n4533 );
not ( n4535 , n2315 );
nand ( n4536 , n4535 , n1006 );
not ( n4537 , n4536 );
not ( n4538 , n4501 );
nand ( n4539 , n4537 , n4538 );
nand ( n4540 , n4534 , n4539 );
nor ( n4541 , n4530 , n4540 );
not ( n4542 , n4541 );
nand ( n4543 , n4542 , n4520 , n4514 , n4521 );
nand ( n4544 , n4518 , n4522 , n4543 );
not ( n4545 , n4544 );
nand ( n4546 , n4505 , n4541 );
not ( n4547 , n4502 );
nand ( n4548 , n1025 , n4453 );
nand ( n4549 , n4548 , n4444 );
not ( n4550 , n4549 );
nand ( n4551 , n4546 , n4547 , n4550 );
not ( n4552 , n4300 );
and ( n4553 , n4552 , n4470 );
not ( n4554 , n4512 );
not ( n4555 , n4554 );
and ( n4556 , n4553 , n4555 , n4516 );
nand ( n4557 , n4556 , n4506 );
not ( n4558 , n26 );
not ( n4559 , n4299 );
and ( n4560 , n4558 , n4512 , n4559 );
nand ( n4561 , n4560 , n4550 );
not ( n4562 , n4560 );
not ( n4563 , n4513 );
not ( n4564 , n4563 );
or ( n4565 , n4562 , n4564 );
not ( n4566 , n26 );
nand ( n4567 , n4566 , n4454 );
nand ( n4568 , n4565 , n4567 );
nand ( n4569 , n4521 , n4568 );
and ( n4570 , n4551 , n4557 , n4561 , n4569 );
nand ( n4571 , n4553 , n4555 , n4516 );
nor ( n4572 , n4571 , n4541 );
nor ( n4573 , n4519 , n4549 );
not ( n4574 , n4573 );
not ( n4575 , n4546 );
or ( n4576 , n4574 , n4575 );
nand ( n4577 , n4576 , n35 );
nor ( n4578 , n4572 , n4577 );
nand ( n4579 , n4545 , n4570 , n4578 );
nand ( n4580 , n4509 , n4579 );
not ( n4581 , n4580 );
or ( n4582 , n4485 , n4581 );
nand ( n4583 , n4582 , n4541 );
not ( n4584 , n4579 );
nor ( n4585 , n4583 , n4584 );
not ( n4586 , n4585 );
not ( n4587 , n4586 );
and ( n4588 , n1223 , n4587 );
not ( n4589 , n4484 );
not ( n4590 , n4488 );
not ( n4591 , n4559 );
and ( n4592 , n199 , n4591 );
not ( n4593 , n4336 );
nor ( n4594 , n4592 , n4593 );
not ( n4595 , n4594 );
not ( n4596 , n4595 );
not ( n4597 , n4394 );
nand ( n4598 , n1152 , n4597 );
nand ( n4599 , n4323 , n4596 , n4598 );
not ( n4600 , n4599 );
or ( n4601 , n4590 , n4600 );
not ( n4602 , n26 );
not ( n4603 , n4385 );
and ( n4604 , n4602 , n4603 , n171 , n391 );
nand ( n4605 , n32 , n4346 );
not ( n4606 , n4352 );
not ( n4607 , n4354 );
and ( n4608 , n4605 , n4606 , n4607 );
not ( n4609 , n4608 );
nand ( n4610 , n1025 , n4374 );
nand ( n4611 , n4609 , n4610 );
not ( n4612 , n4611 );
nand ( n4613 , n4604 , n4612 );
not ( n4614 , n4357 );
not ( n4615 , n4604 );
not ( n4616 , n4300 );
not ( n4617 , n177 );
nand ( n4618 , n391 , n389 , n4617 );
nand ( n4619 , n4616 , n4618 );
nor ( n4620 , n4615 , n4619 );
nand ( n4621 , n4614 , n4620 );
and ( n4622 , n4613 , n35 , n4621 );
not ( n4623 , n26 );
nand ( n4624 , n1053 , n4374 );
nand ( n4625 , n4624 , n4356 );
not ( n4626 , n4625 );
nand ( n4627 , n4394 , n4623 , n4626 );
not ( n4628 , n4365 );
and ( n4629 , n160 , n4628 );
nor ( n4630 , n4629 , n4595 );
not ( n4631 , n4619 );
not ( n4632 , n4357 );
and ( n4633 , n4631 , n4632 );
and ( n4634 , n4630 , n4633 );
not ( n4635 , n4608 );
not ( n4636 , n26 );
and ( n4637 , n4636 , n4346 );
nand ( n4638 , n4635 , n4637 , n4373 );
not ( n4639 , n4638 );
nor ( n4640 , n4634 , n4639 );
and ( n4641 , n4622 , n4627 , n4640 );
not ( n4642 , n4527 );
not ( n4643 , n4365 );
and ( n4644 , n4642 , n4643 );
and ( n4645 , n4537 , n4300 );
nor ( n4646 , n4645 , n4533 );
not ( n4647 , n4646 );
nor ( n4648 , n4644 , n4647 );
not ( n4649 , n4648 );
nor ( n4650 , n4649 , n4630 );
nand ( n4651 , n4375 , n4358 );
not ( n4652 , n4651 );
nor ( n4653 , n4302 , n4611 );
nor ( n4654 , n4652 , n4653 );
nor ( n4655 , n4650 , n4654 );
not ( n4656 , n4366 );
nand ( n4657 , n4656 , n4626 );
or ( n4658 , n4657 , n4650 );
not ( n4659 , n4648 );
nand ( n4660 , n4659 , n4633 );
nand ( n4661 , n4658 , n4660 );
nor ( n4662 , n4655 , n4661 );
nand ( n4663 , n4641 , n4662 );
nand ( n4664 , n4601 , n4663 );
not ( n4665 , n4664 );
or ( n4666 , n4589 , n4665 );
not ( n4667 , n4649 );
nand ( n4668 , n4666 , n4667 );
not ( n4669 , n4663 );
nor ( n4670 , n4668 , n4669 );
not ( n4671 , n4670 );
or ( n4672 , n1913 , n4671 );
nor ( n4673 , n4514 , n4456 );
nor ( n4674 , n4447 , n4673 );
not ( n4675 , n4292 );
nor ( n4676 , n4337 , n4380 );
not ( n4677 , n4676 );
not ( n4678 , n4513 );
not ( n4679 , n4678 );
or ( n4680 , n4677 , n4679 );
nand ( n4681 , n4680 , n4389 );
not ( n4682 , n4681 );
or ( n4683 , n4675 , n4682 );
nand ( n4684 , n4393 , n4497 );
nand ( n4685 , n4683 , n4684 );
nand ( n4686 , n4674 , n4685 );
or ( n4687 , n1143 , n4686 );
nand ( n4688 , n4672 , n4687 );
nor ( n4689 , n4588 , n4688 );
and ( n4690 , n4616 , n4470 );
not ( n4691 , n26 );
nand ( n4692 , n4690 , n4691 , n4516 );
or ( n4693 , n4519 , n4692 );
not ( n4694 , n4526 );
not ( n4695 , n4471 );
or ( n4696 , n4694 , n4695 );
nand ( n4697 , n4696 , n4646 );
not ( n4698 , n4697 );
not ( n4699 , n158 );
not ( n4700 , n4471 );
or ( n4701 , n4699 , n4700 );
nand ( n4702 , n4701 , n4594 );
nand ( n4703 , n4698 , n4702 );
buf ( n4704 , n4548 );
buf ( n4705 , n4704 );
and ( n4706 , n4301 , n4516 );
nand ( n4707 , n4703 , n4705 , n4706 );
not ( n4708 , n4702 );
nand ( n4709 , n4708 , n4515 );
not ( n4710 , n4709 );
nand ( n4711 , n4515 , n4697 );
not ( n4712 , n4711 );
or ( n4713 , n4710 , n4712 );
not ( n4714 , n4445 );
nand ( n4715 , n4461 , n4714 );
not ( n4716 , n4715 );
nand ( n4717 , n4713 , n4716 );
nand ( n4718 , n4693 , n4707 , n4717 );
not ( n4719 , n4718 );
not ( n4720 , n26 );
not ( n4721 , n4453 );
and ( n4722 , n4720 , n4721 , n4516 );
not ( n4723 , n4550 );
not ( n4724 , n4709 );
not ( n4725 , n4724 );
or ( n4726 , n4723 , n4725 );
and ( n4727 , n35 , n4692 );
nand ( n4728 , n4726 , n4727 );
nor ( n4729 , n4722 , n4728 );
or ( n4730 , n4549 , n4711 );
buf ( n4731 , n4603 );
and ( n4732 , n171 , n391 , n4731 , n4470 );
and ( n4733 , n4732 , n4516 );
and ( n4734 , n4733 , n4703 );
not ( n4735 , n4705 );
buf ( n4736 , n4444 );
nand ( n4737 , n4604 , n4736 );
nor ( n4738 , n4735 , n4737 );
nor ( n4739 , n4734 , n4738 );
nand ( n4740 , n4719 , n4729 , n4730 , n4739 );
not ( n4741 , n4488 );
not ( n4742 , n4702 );
nand ( n4743 , n4323 , n4742 );
not ( n4744 , n4743 );
or ( n4745 , n4741 , n4744 );
nand ( n4746 , n4745 , n4740 );
and ( n4747 , n4746 , n4484 );
nor ( n4748 , n4747 , n4697 );
nand ( n4749 , n4740 , n4748 );
not ( n4750 , n4749 );
and ( n4751 , n1909 , n4750 );
not ( n4752 , n4642 );
not ( n4753 , n34 );
not ( n4754 , n4406 );
or ( n4755 , n4753 , n4754 );
not ( n4756 , n4412 );
nand ( n4757 , n4755 , n4756 );
not ( n4758 , n4757 );
not ( n4759 , n4758 );
not ( n4760 , n4759 );
or ( n4761 , n4752 , n4760 );
not ( n4762 , n4534 );
not ( n4763 , n4539 );
nor ( n4764 , n4762 , n4763 );
nand ( n4765 , n4761 , n4764 );
not ( n4766 , n4765 );
not ( n4767 , n4560 );
or ( n4768 , n4767 , n4611 );
not ( n4769 , n4357 );
and ( n4770 , n4560 , n4769 );
nand ( n4771 , n4414 , n4770 );
nand ( n4772 , n4768 , n35 , n4771 );
not ( n4773 , n4758 );
and ( n4774 , n538 , n4773 );
not ( n4775 , n4504 );
nor ( n4776 , n4774 , n4775 );
not ( n4777 , n4776 );
and ( n4778 , n4777 , n4766 );
not ( n4779 , n4651 );
nor ( n4780 , n4502 , n4611 );
nor ( n4781 , n4779 , n4780 );
nor ( n4782 , n4778 , n4781 );
nor ( n4783 , n4772 , n4782 );
not ( n4784 , n4773 );
not ( n4785 , n26 );
nand ( n4786 , n4785 , n4626 );
not ( n4787 , n4786 );
and ( n4788 , n4784 , n4787 );
nor ( n4789 , n4788 , n4639 );
not ( n4790 , n4616 );
nor ( n4791 , n4554 , n4790 );
nand ( n4792 , n4791 , n4614 , n4413 );
not ( n4793 , n4792 );
nand ( n4794 , n4793 , n4765 );
nand ( n4795 , n4789 , n4794 );
nand ( n4796 , n4414 , n4626 );
not ( n4797 , n4796 );
nand ( n4798 , n4765 , n4797 );
not ( n4799 , n4792 );
not ( n4800 , n4796 );
or ( n4801 , n4799 , n4800 );
nand ( n4802 , n4801 , n4776 );
nand ( n4803 , n4798 , n4802 );
nor ( n4804 , n4795 , n4803 );
nand ( n4805 , n4783 , n4804 );
nand ( n4806 , n4766 , n4805 );
not ( n4807 , n4806 );
not ( n4808 , n4488 );
not ( n4809 , n4777 );
nand ( n4810 , n4323 , n4809 );
not ( n4811 , n4810 );
or ( n4812 , n4808 , n4811 );
nand ( n4813 , n4812 , n4805 );
nand ( n4814 , n4484 , n4813 );
nand ( n4815 , n4807 , n4814 );
not ( n4816 , n4815 );
and ( n4817 , n1137 , n4816 );
not ( n4818 , n1880 );
not ( n4819 , n35 );
nand ( n4820 , n4819 , n4487 );
not ( n4821 , n4820 );
and ( n4822 , n158 , n4538 );
nor ( n4823 , n4822 , n4337 );
buf ( n4824 , n4823 );
not ( n4825 , n4495 );
not ( n4826 , n200 );
nand ( n4827 , n4825 , n4826 );
nand ( n4828 , n4824 , n4322 , n4827 );
not ( n4829 , n4828 );
or ( n4830 , n4821 , n4829 );
not ( n4831 , n4537 );
not ( n4832 , n4496 );
or ( n4833 , n4831 , n4832 );
and ( n4834 , n4526 , n4502 );
nor ( n4835 , n4834 , n4533 );
nand ( n4836 , n4833 , n4835 );
not ( n4837 , n4836 );
and ( n4838 , n4704 , n4678 , n4736 );
not ( n4839 , n4838 );
or ( n4840 , n4837 , n4839 );
not ( n4841 , n26 );
nand ( n4842 , n4841 , n4714 , n4704 , n4678 );
nand ( n4843 , n4840 , n4842 );
nand ( n4844 , n4823 , n4827 );
not ( n4845 , n4844 );
not ( n4846 , n4845 );
not ( n4847 , n4838 );
or ( n4848 , n4846 , n4847 );
not ( n4849 , n4836 );
nand ( n4850 , n4844 , n4849 );
not ( n4851 , n4555 );
nor ( n4852 , n4851 , n4302 );
nand ( n4853 , n4850 , n4517 , n4852 );
nand ( n4854 , n4848 , n4853 );
nor ( n4855 , n4843 , n4854 );
nand ( n4856 , n4824 , n4827 , n4556 );
nand ( n4857 , n4560 , n4517 );
nand ( n4858 , n4856 , n4857 , n4569 );
nor ( n4859 , n4571 , n4849 );
not ( n4860 , n4859 );
not ( n4861 , n35 );
not ( n4862 , n4515 );
nor ( n4863 , n4862 , n4549 );
not ( n4864 , n4823 );
not ( n4865 , n4827 );
or ( n4866 , n4864 , n4865 );
nand ( n4867 , n4866 , n4849 );
nand ( n4868 , n4863 , n4867 );
nand ( n4869 , n4860 , n4861 , n4868 );
nor ( n4870 , n4858 , n4869 );
nand ( n4871 , n4855 , n4870 );
nand ( n4872 , n4830 , n4871 );
and ( n4873 , n4872 , n4484 );
not ( n4874 , n4871 );
nor ( n4875 , n4873 , n4874 );
nand ( n4876 , n4875 , n4849 );
not ( n4877 , n4876 );
and ( n4878 , n4818 , n4877 );
not ( n4879 , n19 );
not ( n4880 , n23 );
nor ( n4881 , n4879 , n4880 );
nor ( n4882 , n4878 , n4881 );
not ( n4883 , n1375 );
nand ( n4884 , n4322 , n1382 , n4547 );
buf ( n4885 , n4731 );
and ( n4886 , n234 , n4314 );
nand ( n4887 , n171 , n4885 , n4886 );
not ( n4888 , n4554 );
nand ( n4889 , n4888 , n4314 , n4465 , n4301 );
nand ( n4890 , n4887 , n4889 );
nand ( n4891 , n4292 , n4890 );
and ( n4892 , n4884 , n4891 );
not ( n4893 , n4892 );
and ( n4894 , n4883 , n4893 );
nand ( n4895 , n4560 , n4626 );
not ( n4896 , n35 );
and ( n4897 , n4895 , n4896 , n4771 );
not ( n4898 , n201 );
not ( n4899 , n4757 );
or ( n4900 , n4898 , n4899 );
nand ( n4901 , n4900 , n4824 );
not ( n4902 , n4901 );
and ( n4903 , n4902 , n4793 );
not ( n4904 , n4414 );
nor ( n4905 , n4611 , n26 );
not ( n4906 , n4905 );
or ( n4907 , n4904 , n4906 );
nand ( n4908 , n4907 , n4638 );
nor ( n4909 , n4903 , n4908 );
nand ( n4910 , n4897 , n4909 );
not ( n4911 , n4537 );
not ( n4912 , n4757 );
or ( n4913 , n4911 , n4912 );
nor ( n4914 , n4525 , n4501 );
nor ( n4915 , n4762 , n4914 );
nand ( n4916 , n4913 , n4915 );
not ( n4917 , n4916 );
nand ( n4918 , n4901 , n4917 );
nor ( n4919 , n4851 , n4302 );
nand ( n4920 , n4918 , n4626 , n4919 );
nand ( n4921 , n4793 , n4916 );
not ( n4922 , n4651 );
nand ( n4923 , n4414 , n4610 , n4358 );
not ( n4924 , n4923 );
or ( n4925 , n4922 , n4924 );
nand ( n4926 , n4925 , n4918 );
nand ( n4927 , n4920 , n4921 , n4926 );
or ( n4928 , n4910 , n4927 );
not ( n4929 , n534 );
or ( n4930 , n4929 , n4414 );
nand ( n4931 , n4930 , n4322 , n4824 );
nand ( n4932 , n4820 , n4931 );
nand ( n4933 , n4928 , n4932 );
and ( n4934 , n4933 , n4484 );
or ( n4935 , n4910 , n4927 );
nand ( n4936 , n4935 , n4917 );
nor ( n4937 , n4934 , n4936 );
and ( n4938 , n764 , n4937 );
nor ( n4939 , n4894 , n4938 );
nand ( n4940 , n4882 , n4939 );
not ( n4941 , n4940 );
or ( n4942 , n1371 , n4941 );
nand ( n4943 , n4394 , n4905 );
nand ( n4944 , n4826 , n4619 );
not ( n4945 , n4559 );
nand ( n4946 , n158 , n4945 );
nand ( n4947 , n4944 , n4465 , n4946 );
not ( n4948 , n4947 );
nand ( n4949 , n4948 , n4633 );
nand ( n4950 , n4943 , n4638 , n4949 );
not ( n4951 , n4950 );
not ( n4952 , n4365 );
and ( n4953 , n4537 , n4952 );
not ( n4954 , n4525 );
not ( n4955 , n4559 );
and ( n4956 , n4954 , n4955 );
nor ( n4957 , n4956 , n4533 );
not ( n4958 , n4957 );
nor ( n4959 , n4953 , n4958 );
nand ( n4960 , n4947 , n4959 );
not ( n4961 , n4358 );
and ( n4962 , n4631 , n4610 );
not ( n4963 , n4962 );
or ( n4964 , n4961 , n4963 );
nand ( n4965 , n4964 , n4651 );
and ( n4966 , n4960 , n4965 );
not ( n4967 , n4604 );
not ( n4968 , n4626 );
or ( n4969 , n4967 , n4968 );
not ( n4970 , n4621 );
nor ( n4971 , n35 , n4970 );
nand ( n4972 , n4969 , n4971 );
nor ( n4973 , n4966 , n4972 );
not ( n4974 , n4959 );
nand ( n4975 , n4633 , n4974 );
not ( n4976 , n4624 );
nor ( n4977 , n4302 , n4976 );
nand ( n4978 , n4977 , n4358 , n4960 );
nand ( n4979 , n4951 , n4973 , n4975 , n4978 );
not ( n4980 , n4820 );
nand ( n4981 , n4465 , n4946 );
not ( n4982 , n4981 );
nand ( n4983 , n4322 , n4982 , n4944 );
not ( n4984 , n4983 );
or ( n4985 , n4980 , n4984 );
nand ( n4986 , n4985 , n4979 );
and ( n4987 , n4484 , n4986 );
nor ( n4988 , n4987 , n4974 );
nand ( n4989 , n4979 , n4988 );
not ( n4990 , n4989 );
and ( n4991 , n590 , n4990 );
nand ( n4992 , n4826 , n4471 );
nand ( n4993 , n4315 , n4982 , n4992 );
nand ( n4994 , n4820 , n4993 );
not ( n4995 , n4994 );
and ( n4996 , n4484 , n4995 );
not ( n4997 , n4537 );
not ( n4998 , n4471 );
or ( n4999 , n4997 , n4998 );
nand ( n5000 , n4999 , n4957 );
nor ( n5001 , n4996 , n5000 );
not ( n5002 , n35 );
nand ( n5003 , n4732 , n4714 , n4982 , n4992 );
and ( n5004 , n4733 , n5000 );
not ( n5005 , n4704 );
nor ( n5006 , n5005 , n4692 );
nor ( n5007 , n5004 , n5006 );
and ( n5008 , n5002 , n4692 , n5003 , n5007 );
nand ( n5009 , n4982 , n4992 , n4454 , n4736 );
not ( n5010 , n4722 );
nand ( n5011 , n4714 , n4454 , n5000 );
nand ( n5012 , n5009 , n5010 , n5011 );
not ( n5013 , n4520 );
not ( n5014 , n4981 );
not ( n5015 , n5014 );
not ( n5016 , n4992 );
or ( n5017 , n5015 , n5016 );
not ( n5018 , n5000 );
nand ( n5019 , n5017 , n5018 );
and ( n5020 , n4706 , n5019 );
not ( n5021 , n4737 );
nor ( n5022 , n5020 , n5021 );
or ( n5023 , n5013 , n5022 );
not ( n5024 , n4715 );
nand ( n5025 , n5024 , n5019 , n4705 );
nand ( n5026 , n5023 , n5025 );
nor ( n5027 , n5012 , n5026 );
nand ( n5028 , n5008 , n5027 );
and ( n5029 , n5001 , n5028 );
not ( n5030 , n5029 );
or ( n5031 , n521 , n5030 );
not ( n5032 , n16 );
nand ( n5033 , n23 , n5032 );
nand ( n5034 , n5031 , n5033 );
nor ( n5035 , n4991 , n5034 );
or ( n5036 , n1415 , n5035 );
nand ( n5037 , n4942 , n5036 );
nor ( n5038 , n4751 , n4817 , n5037 );
and ( n5039 , n4483 , n4689 , n5038 );
nor ( n5040 , n5039 , n1971 );
not ( n5041 , n1849 );
not ( n5042 , n21 );
not ( n5043 , n24 );
and ( n5044 , n2316 , n4406 );
not ( n5045 , n2316 );
not ( n5046 , n4306 );
and ( n5047 , n5045 , n5046 );
nor ( n5048 , n5044 , n5047 );
not ( n5049 , n5048 );
nand ( n5050 , n5043 , n5049 );
or ( n5051 , n5042 , n5050 );
not ( n5052 , n5051 );
not ( n5053 , n5052 );
not ( n5054 , n5053 );
not ( n5055 , n5054 );
not ( n5056 , n5055 );
not ( n5057 , n4876 );
not ( n5058 , n5057 );
or ( n5059 , n5056 , n5058 );
not ( n5060 , n23 );
nor ( n5061 , n22 , n24 );
not ( n5062 , n21 );
nor ( n5063 , n5062 , n31 );
nand ( n5064 , n5050 , n5061 , n5063 );
nand ( n5065 , n5060 , n5064 );
not ( n5066 , n5065 );
buf ( n5067 , n5066 );
buf ( n5068 , n5067 );
buf ( n5069 , n5068 );
nand ( n5070 , n5059 , n5069 );
and ( n5071 , n5070 , n1432 );
not ( n5072 , n5051 );
not ( n5073 , n5072 );
not ( n5074 , n5073 );
not ( n5075 , n4427 );
or ( n5076 , n5074 , n5075 );
nand ( n5077 , n5076 , n5067 );
and ( n5078 , n1613 , n5077 );
nor ( n5079 , n5071 , n5078 );
not ( n5080 , n5053 );
not ( n5081 , n5080 );
not ( n5082 , n4580 );
nand ( n5083 , n5081 , n5082 );
nand ( n5084 , n5068 , n5083 );
and ( n5085 , n1559 , n5084 );
not ( n5086 , n1556 );
or ( n5087 , n5054 , n4746 );
not ( n5088 , n5067 );
not ( n5089 , n5088 );
nand ( n5090 , n5087 , n5089 );
not ( n5091 , n5090 );
or ( n5092 , n5086 , n5091 );
not ( n5093 , n5028 );
or ( n5094 , n5093 , n5052 , n4995 );
nand ( n5095 , n5094 , n5066 );
nand ( n5096 , n1621 , n5095 );
nand ( n5097 , n5092 , n5096 );
or ( n5098 , n5080 , n4933 );
nand ( n5099 , n5098 , n5089 );
not ( n5100 , n5099 );
nor ( n5101 , n1572 , n5100 );
nor ( n5102 , n5085 , n5097 , n5101 );
nand ( n5103 , n17 , n692 );
nand ( n5104 , n23 , n5103 );
or ( n5105 , n1371 , n5104 );
not ( n5106 , n5073 );
not ( n5107 , n4886 );
or ( n5108 , n4307 , n5107 );
nand ( n5109 , n5108 , n4889 );
not ( n5110 , n5109 );
or ( n5111 , n5106 , n5110 );
nand ( n5112 , n5111 , n5067 );
and ( n5113 , n1590 , n5112 );
and ( n5114 , n114 , n5049 );
or ( n5115 , n4318 , n5114 );
not ( n5116 , n5065 );
nand ( n5117 , n5115 , n5116 );
and ( n5118 , n1592 , n5117 );
nor ( n5119 , n5113 , n5118 );
not ( n5120 , n18 );
not ( n5121 , n1589 );
not ( n5122 , n5073 );
or ( n5123 , n5122 , n4892 );
nand ( n5124 , n5123 , n5067 );
nand ( n5125 , n5120 , n5121 , n5124 );
nand ( n5126 , n5105 , n5119 , n5125 );
and ( n5127 , n16 , n1314 );
not ( n5128 , n1409 );
nor ( n5129 , n5127 , n5128 , n1416 );
or ( n5130 , n5104 , n5129 );
not ( n5131 , n1550 );
and ( n5132 , n4423 , n5051 , n4416 );
nor ( n5133 , n5132 , n5065 );
or ( n5134 , n5131 , n5133 );
and ( n5135 , n4674 , n5051 , n4681 );
nor ( n5136 , n5135 , n5065 );
or ( n5137 , n1563 , n5136 );
nand ( n5138 , n5130 , n5134 , n5137 );
nor ( n5139 , n5126 , n5138 );
not ( n5140 , n5122 );
not ( n5141 , n4813 );
nand ( n5142 , n5140 , n5141 );
nand ( n5143 , n5068 , n5142 );
not ( n5144 , n5143 );
or ( n5145 , n5144 , n1542 );
not ( n5146 , n308 );
not ( n5147 , n1583 );
or ( n5148 , n5146 , n5147 );
not ( n5149 , n5104 );
nand ( n5150 , n5148 , n5149 );
not ( n5151 , n4986 );
not ( n5152 , n5151 );
or ( n5153 , n5122 , n5152 );
nand ( n5154 , n5153 , n5067 );
nand ( n5155 , n1623 , n5154 );
nand ( n5156 , n5145 , n5150 , n5155 );
or ( n5157 , n4872 , n5080 );
nand ( n5158 , n5157 , n5067 );
not ( n5159 , n5158 );
or ( n5160 , n1568 , n5159 );
not ( n5161 , n4664 );
nand ( n5162 , n5140 , n5161 );
nand ( n5163 , n5089 , n5162 );
nand ( n5164 , n1627 , n5163 );
buf ( n5165 , n1936 );
not ( n5166 , n5165 );
not ( n5167 , n4378 );
and ( n5168 , n5167 , n5051 , n4390 );
nor ( n5169 , n5168 , n5065 );
or ( n5170 , n5166 , n5169 );
nor ( n5171 , n4447 , n4462 );
and ( n5172 , n5171 , n5051 , n4473 );
nor ( n5173 , n5172 , n5065 );
or ( n5174 , n795 , n5173 );
nand ( n5175 , n5170 , n5174 );
and ( n5176 , n1582 , n5175 );
or ( n5177 , n16 , n1575 );
not ( n5178 , n1600 );
nand ( n5179 , n5177 , n5178 );
and ( n5180 , n5149 , n5179 );
nor ( n5181 , n5176 , n5180 );
nand ( n5182 , n5160 , n5164 , n5181 );
nor ( n5183 , n5156 , n5182 );
and ( n5184 , n5079 , n5102 , n5139 , n5183 );
nand ( n5185 , n5055 , n4585 );
nand ( n5186 , n5069 , n5185 );
and ( n5187 , n5186 , n1223 );
not ( n5188 , n5055 );
not ( n5189 , n4750 );
or ( n5190 , n5188 , n5189 );
nand ( n5191 , n5190 , n5069 );
and ( n5192 , n1317 , n5191 );
nor ( n5193 , n5187 , n5192 );
or ( n5194 , n5052 , n4397 );
nand ( n5195 , n5194 , n5066 );
and ( n5196 , n14 , n5195 );
not ( n5197 , n14 );
or ( n5198 , n5052 , n4479 );
nand ( n5199 , n5198 , n5066 );
and ( n5200 , n5197 , n5199 );
nor ( n5201 , n5196 , n5200 );
nor ( n5202 , n432 , n5201 );
and ( n5203 , n1406 , n5202 );
not ( n5204 , n5053 );
not ( n5205 , n4326 );
or ( n5206 , n5204 , n5205 );
nand ( n5207 , n5206 , n5067 );
and ( n5208 , n1419 , n5207 );
nor ( n5209 , n5203 , n5208 );
not ( n5210 , n5054 );
not ( n5211 , n5210 );
not ( n5212 , n4990 );
or ( n5213 , n5211 , n5212 );
nand ( n5214 , n5213 , n5069 );
and ( n5215 , n1837 , n5214 );
nand ( n5216 , n5055 , n4670 );
nand ( n5217 , n5216 , n5069 );
and ( n5218 , n5217 , n1319 );
nor ( n5219 , n5215 , n5218 );
and ( n5220 , n5209 , n5219 );
nand ( n5221 , n5210 , n4816 );
nand ( n5222 , n5069 , n5221 );
and ( n5223 , n1137 , n5222 );
or ( n5224 , n5072 , n4686 );
nand ( n5225 , n5224 , n5066 );
and ( n5226 , n1144 , n5225 );
not ( n5227 , n5029 );
or ( n5228 , n5227 , n5080 );
not ( n5229 , n5088 );
nand ( n5230 , n5228 , n5229 );
nand ( n5231 , n5230 , n1730 , n520 );
not ( n5232 , n5210 );
not ( n5233 , n4937 );
or ( n5234 , n5232 , n5233 );
nand ( n5235 , n5234 , n5069 );
nand ( n5236 , n1787 , n5235 );
nand ( n5237 , n5231 , n5236 );
nor ( n5238 , n5223 , n5226 , n5237 );
nand ( n5239 , n5184 , n5193 , n5220 , n5238 );
not ( n5240 , n5239 );
or ( n5241 , n5041 , n5240 );
not ( n5242 , n5141 );
not ( n5243 , n5242 );
not ( n5244 , n5243 );
or ( n5245 , n2011 , n5244 );
nand ( n5246 , n5241 , n5245 );
nor ( n5247 , n5040 , n5246 );
not ( n5248 , n5082 );
not ( n5249 , n5248 );
and ( n5250 , n2028 , n5249 );
not ( n5251 , n23 );
or ( n5252 , n5251 , n1971 , n1583 );
not ( n5253 , n4473 );
not ( n5254 , n5253 );
nand ( n5255 , n5171 , n2023 , n5254 );
nand ( n5256 , n5252 , n5255 );
not ( n5257 , n4417 );
not ( n5258 , n5257 );
not ( n5259 , n5258 );
and ( n5260 , n4423 , n2018 , n5259 );
nor ( n5261 , n5250 , n5256 , n5260 );
not ( n5262 , n4933 );
and ( n5263 , n764 , n5262 );
nor ( n5264 , n5263 , n4881 );
buf ( n5265 , n4872 );
not ( n5266 , n5265 );
and ( n5267 , n583 , n5266 );
and ( n5268 , n1374 , n4890 );
nor ( n5269 , n5267 , n5268 );
nand ( n5270 , n5264 , n5269 );
and ( n5271 , n2033 , n5270 );
and ( n5272 , n590 , n5151 );
nor ( n5273 , n5093 , n521 , n4995 );
not ( n5274 , n5033 );
nor ( n5275 , n5272 , n5273 , n5274 );
not ( n5276 , n5275 );
and ( n5277 , n2041 , n5276 );
nor ( n5278 , n5271 , n5277 );
not ( n5279 , n5161 );
not ( n5280 , n5279 );
and ( n5281 , n2030 , n5280 );
not ( n5282 , n4746 );
and ( n5283 , n2014 , n5282 );
not ( n5284 , n4674 );
not ( n5285 , n5284 );
not ( n5286 , n4681 );
not ( n5287 , n5286 );
not ( n5288 , n5287 );
not ( n5289 , n5288 );
and ( n5290 , n5285 , n1998 , n5289 );
not ( n5291 , n4390 );
not ( n5292 , n5291 );
not ( n5293 , n5292 );
not ( n5294 , n5293 );
and ( n5295 , n5167 , n2004 , n5294 );
nor ( n5296 , n5290 , n5295 );
not ( n5297 , n5296 );
nor ( n5298 , n5281 , n5283 , n5297 );
not ( n5299 , n1990 );
not ( n5300 , n4318 );
and ( n5301 , n5299 , n5300 );
and ( n5302 , n4330 , n2010 );
nor ( n5303 , n5301 , n5302 );
nand ( n5304 , n23 , n1852 , n1600 );
nand ( n5305 , n18 , n23 , n1852 , n3256 );
and ( n5306 , n5298 , n5303 , n5304 , n5305 );
nand ( n5307 , n5247 , n5261 , n5278 , n5306 );
not ( n5308 , n5307 );
not ( n5309 , n5308 );
and ( n5310 , n4280 , n5309 );
and ( n5311 , n2618 , n5084 );
not ( n5312 , n313 );
not ( n5313 , n5312 );
not ( n5314 , n5313 );
not ( n5315 , n5314 );
not ( n5316 , n5315 );
not ( n5317 , n5316 );
or ( n5318 , n5166 , n5133 );
or ( n5319 , n795 , n5136 );
nand ( n5320 , n5318 , n5319 );
and ( n5321 , n5317 , n5320 );
nor ( n5322 , n795 , n5114 );
nand ( n5323 , n5285 , n5322 , n5287 );
not ( n5324 , n5165 );
nor ( n5325 , n5324 , n5114 );
nand ( n5326 , n4423 , n5325 , n5257 );
nand ( n5327 , n5323 , n5326 );
not ( n5328 , n312 );
not ( n5329 , n5328 );
not ( n5330 , n5329 );
not ( n5331 , n5330 );
nor ( n5332 , n5331 , n1995 );
nor ( n5333 , n5321 , n5327 , n5332 );
not ( n5334 , n5333 );
and ( n5335 , n2726 , n5334 );
nor ( n5336 , n5311 , n5335 );
not ( n5337 , n766 );
not ( n5338 , n5099 );
or ( n5339 , n5337 , n5338 );
and ( n5340 , n5158 , n584 );
and ( n5341 , n782 , n5112 );
nor ( n5342 , n5340 , n5341 );
nand ( n5343 , n5339 , n5342 );
and ( n5344 , n2582 , n5343 );
not ( n5345 , n5316 );
not ( n5346 , n5345 );
buf ( n5347 , n5346 );
not ( n5348 , n5347 );
and ( n5349 , n5348 , n5084 );
not ( n5350 , n5331 );
not ( n5351 , n5350 );
not ( n5352 , n5351 );
not ( n5353 , n5352 );
nand ( n5354 , n5353 , n5083 );
nor ( n5355 , n5349 , n5354 );
nor ( n5356 , n5355 , n2604 , n2624 );
nor ( n5357 , n5344 , n5356 );
nand ( n5358 , n5336 , n5357 );
nor ( n5359 , n765 , n5114 );
and ( n5360 , n5359 , n5262 );
not ( n5361 , n5114 );
nand ( n5362 , n584 , n5361 );
or ( n5363 , n5362 , n5265 );
not ( n5364 , n5210 );
nand ( n5365 , n570 , n4890 );
or ( n5366 , n5364 , n5365 );
nand ( n5367 , n5330 , n520 );
not ( n5368 , n633 );
nand ( n5369 , n5330 , n5368 );
and ( n5370 , n5367 , n5369 );
nor ( n5371 , n5370 , n625 );
not ( n5372 , n5371 );
nand ( n5373 , n5363 , n5366 , n5372 );
nor ( n5374 , n5360 , n5373 );
not ( n5375 , n5346 );
nand ( n5376 , n5375 , n5343 );
and ( n5377 , n5374 , n5376 );
or ( n5378 , n2700 , n5377 );
or ( n5379 , n2583 , n5144 );
nand ( n5380 , n5378 , n5379 );
not ( n5381 , n994 );
not ( n5382 , n5239 );
or ( n5383 , n5381 , n5382 );
and ( n5384 , n5345 , n5143 );
nand ( n5385 , n5351 , n5142 );
nor ( n5386 , n5384 , n5385 );
or ( n5387 , n2588 , n5386 );
nand ( n5388 , n5383 , n5387 );
nor ( n5389 , n5358 , n5380 , n5388 );
nand ( n5390 , n856 , n989 );
or ( n5391 , n5390 , n5333 );
nor ( n5392 , n308 , n3369 );
not ( n5393 , n40 );
nand ( n5394 , n97 , n5392 , n5393 , n5143 );
nand ( n5395 , n5391 , n5394 );
not ( n5396 , n40 );
and ( n5397 , n2615 , n5392 , n5396 , n5084 );
not ( n5398 , n5392 );
not ( n5399 , n40 );
nor ( n5400 , n5398 , n5399 , n5355 , n2616 );
nor ( n5401 , n5395 , n5397 , n5400 );
not ( n5402 , n40 );
and ( n5403 , n5402 , n989 , n5343 );
not ( n5404 , n20 );
not ( n5405 , n5103 );
not ( n5406 , n40 );
not ( n5407 , n298 );
or ( n5408 , n5406 , n5407 );
nand ( n5409 , n5408 , n23 );
nor ( n5410 , n5405 , n5409 );
nand ( n5411 , n5404 , n5410 );
nor ( n5412 , n3440 , n5411 );
nor ( n5413 , n5403 , n5412 );
and ( n5414 , n5320 , n853 , n989 );
not ( n5415 , n914 );
not ( n5416 , n5154 );
or ( n5417 , n5415 , n5416 );
and ( n5418 , n909 , n5095 );
and ( n5419 , n942 , n5117 );
nor ( n5420 , n5418 , n5419 );
nand ( n5421 , n5417 , n5420 );
and ( n5422 , n287 , n5421 );
not ( n5423 , n83 );
not ( n5424 , n311 );
or ( n5425 , n5423 , n5424 );
not ( n5426 , n23 );
not ( n5427 , n84 );
or ( n5428 , n5426 , n5427 );
nand ( n5429 , n5425 , n5428 );
not ( n5430 , n5429 );
nor ( n5431 , n5430 , n5405 , n2600 );
and ( n5432 , n20 , n5431 );
nand ( n5433 , n14 , n5103 );
or ( n5434 , n2067 , n5433 , n5430 );
or ( n5435 , n5430 , n912 , n5405 );
nand ( n5436 , n5434 , n5435 );
nor ( n5437 , n5422 , n5432 , n5436 );
and ( n5438 , n5375 , n5163 );
not ( n5439 , n5353 );
not ( n5440 , n5162 );
nor ( n5441 , n5438 , n5439 , n5440 );
not ( n5442 , n5441 );
not ( n5443 , n2653 );
nor ( n5444 , n41 , n5443 );
nand ( n5445 , n5442 , n5444 );
nor ( n5446 , n2616 , n5114 );
and ( n5447 , n5446 , n5282 );
not ( n5448 , n5291 );
and ( n5449 , n5167 , n5325 , n5448 );
or ( n5450 , n5332 , n5449 );
nor ( n5451 , n5447 , n5450 );
nor ( n5452 , n5316 , n2616 );
and ( n5453 , n5452 , n5090 );
not ( n5454 , n5175 );
or ( n5455 , n5316 , n5454 );
nand ( n5456 , n5350 , n2615 );
nand ( n5457 , n5455 , n5456 );
and ( n5458 , n5171 , n5322 , n5254 );
nor ( n5459 , n5453 , n5457 , n5458 );
nand ( n5460 , n5451 , n5459 );
and ( n5461 , n2077 , n5460 );
not ( n5462 , n2615 );
not ( n5463 , n5090 );
or ( n5464 , n5462 , n5463 );
nand ( n5465 , n5464 , n5454 );
and ( n5466 , n2074 , n5465 );
nor ( n5467 , n5461 , n5466 );
nand ( n5468 , n908 , n5350 );
nor ( n5469 , n5468 , n633 );
nand ( n5470 , n909 , n5361 );
or ( n5471 , n5093 , n5470 , n4995 );
or ( n5472 , n4318 , n963 , n5054 );
nand ( n5473 , n5471 , n5472 );
nor ( n5474 , n5469 , n5473 );
not ( n5475 , n912 );
not ( n5476 , n5367 );
and ( n5477 , n5475 , n5476 );
not ( n5478 , n5345 );
not ( n5479 , n5421 );
or ( n5480 , n5478 , n5479 );
nor ( n5481 , n913 , n5114 );
not ( n5482 , n5152 );
nand ( n5483 , n5481 , n5482 );
nand ( n5484 , n5480 , n5483 );
nor ( n5485 , n5477 , n5484 );
and ( n5486 , n5474 , n5485 );
nor ( n5487 , n5486 , n40 );
and ( n5488 , n445 , n5487 );
nor ( n5489 , n286 , n2629 );
and ( n5490 , n5489 , n5163 );
nor ( n5491 , n5488 , n5490 );
nand ( n5492 , n5437 , n5445 , n5467 , n5491 );
and ( n5493 , n442 , n5492 );
nor ( n5494 , n5414 , n5493 );
and ( n5495 , n5389 , n5401 , n5413 , n5494 );
not ( n5496 , n40 );
or ( n5497 , n5496 , n3440 , n5377 );
nand ( n5498 , n97 , n5392 );
not ( n5499 , n40 );
or ( n5500 , n5498 , n5499 , n5386 );
nand ( n5501 , n5497 , n5500 );
not ( n5502 , n5501 );
nor ( n5503 , n5432 , n5436 );
not ( n5504 , n5191 );
or ( n5505 , n2616 , n5504 );
not ( n5506 , n5202 );
nand ( n5507 , n5505 , n5506 );
and ( n5508 , n20 , n5507 );
not ( n5509 , n914 );
not ( n5510 , n5214 );
or ( n5511 , n5509 , n5510 );
and ( n5512 , n909 , n5230 );
and ( n5513 , n942 , n5207 );
nor ( n5514 , n5512 , n5513 );
nand ( n5515 , n5511 , n5514 );
nor ( n5516 , n5508 , n5515 );
or ( n5517 , n2056 , n5516 );
not ( n5518 , n5347 );
and ( n5519 , n5518 , n5217 );
not ( n5520 , n5439 );
nand ( n5521 , n5520 , n5216 );
nor ( n5522 , n5519 , n5521 );
not ( n5523 , n5522 );
and ( n5524 , n5444 , n5523 );
and ( n5525 , n5489 , n5217 );
nor ( n5526 , n5524 , n5525 );
not ( n5527 , n40 );
and ( n5528 , n5481 , n4990 );
nor ( n5529 , n5528 , n5469 );
or ( n5530 , n521 , n5468 );
and ( n5531 , n5361 , n942 , n4326 );
not ( n5532 , n5470 );
not ( n5533 , n5030 );
and ( n5534 , n5532 , n5533 );
nor ( n5535 , n5531 , n5534 );
not ( n5536 , n5347 );
nand ( n5537 , n5536 , n5515 );
nand ( n5538 , n5529 , n5530 , n5535 , n5537 );
and ( n5539 , n5527 , n5538 );
and ( n5540 , n5539 , n445 );
and ( n5541 , n5446 , n4750 );
nor ( n5542 , n5541 , n5332 );
nand ( n5543 , n5322 , n4480 );
and ( n5544 , n5375 , n5202 );
and ( n5545 , n5325 , n4398 );
nor ( n5546 , n5544 , n5545 );
nand ( n5547 , n5452 , n5191 );
and ( n5548 , n5546 , n5456 , n5547 );
and ( n5549 , n5542 , n5543 , n5548 );
not ( n5550 , n5549 );
and ( n5551 , n5550 , n2077 );
nor ( n5552 , n5540 , n5551 );
nand ( n5553 , n5503 , n5517 , n5526 , n5552 );
and ( n5554 , n2121 , n5553 );
not ( n5555 , n442 );
or ( n5556 , n457 , n5355 );
not ( n5557 , n2199 );
not ( n5558 , n5333 );
and ( n5559 , n5557 , n5558 );
and ( n5560 , n511 , n5084 );
nor ( n5561 , n5559 , n5560 );
nand ( n5562 , n5556 , n5561 );
not ( n5563 , n5562 );
not ( n5564 , n20 );
and ( n5565 , n5564 , n99 , n5143 );
or ( n5566 , n20 , n2102 , n5386 );
or ( n5567 , n5377 , n2064 );
nand ( n5568 , n5566 , n5567 );
nor ( n5569 , n5565 , n5568 );
and ( n5570 , n287 , n5343 );
nand ( n5571 , n92 , n5429 );
nor ( n5572 , n2346 , n5571 );
and ( n5573 , n454 , n5572 );
not ( n5574 , n17 );
and ( n5575 , n5574 , n5429 );
and ( n5576 , n2679 , n5575 );
nor ( n5577 , n5570 , n5573 , n5576 );
and ( n5578 , n440 , n5320 );
nor ( n5579 , n5430 , n5405 , n2681 );
not ( n5580 , n3175 );
nor ( n5581 , n5430 , n5580 , n5405 );
nor ( n5582 , n5578 , n5579 , n5581 );
nand ( n5583 , n5563 , n5569 , n5577 , n5582 );
not ( n5584 , n5583 );
or ( n5585 , n5555 , n5584 );
not ( n5586 , n5465 );
or ( n5587 , n868 , n5586 );
not ( n5588 , n40 );
or ( n5589 , n5588 , n5486 );
nand ( n5590 , n20 , n5410 );
nand ( n5591 , n5587 , n5589 , n5590 );
not ( n5592 , n717 );
not ( n5593 , n5441 );
and ( n5594 , n5592 , n5593 );
and ( n5595 , n648 , n5163 );
nor ( n5596 , n5594 , n5595 );
and ( n5597 , n2283 , n5460 );
not ( n5598 , n40 );
and ( n5599 , n5598 , n5421 );
nor ( n5600 , n5597 , n5599 );
nand ( n5601 , n5596 , n5600 );
or ( n5602 , n5591 , n5601 );
nand ( n5603 , n5602 , n989 );
nand ( n5604 , n5585 , n5603 );
nor ( n5605 , n5554 , n5604 );
nand ( n5606 , n5502 , n5605 );
and ( n5607 , n648 , n5217 );
not ( n5608 , n5538 );
not ( n5609 , n40 );
or ( n5610 , n5608 , n5609 );
or ( n5611 , n40 , n5516 );
or ( n5612 , n794 , n5549 );
nand ( n5613 , n5610 , n5611 , n5612 );
or ( n5614 , n717 , n5522 );
nand ( n5615 , n5614 , n5590 );
nor ( n5616 , n5607 , n5613 , n5615 );
or ( n5617 , n2182 , n5616 );
not ( n5618 , n14 );
not ( n5619 , n5618 );
not ( n5620 , n5077 );
and ( n5621 , n5619 , n5620 );
or ( n5622 , n14 , n5225 );
nand ( n5623 , n5622 , n1996 );
nor ( n5624 , n5621 , n5623 );
and ( n5625 , n853 , n5624 );
not ( n5626 , n838 );
and ( n5627 , n5518 , n5186 );
nand ( n5628 , n5520 , n5185 );
nor ( n5629 , n5627 , n5628 );
or ( n5630 , n5626 , n5629 );
nand ( n5631 , n584 , n5070 );
and ( n5632 , n1571 , n5235 );
and ( n5633 , n782 , n5124 );
nor ( n5634 , n5632 , n5633 );
and ( n5635 , n5631 , n5634 );
not ( n5636 , n5635 );
not ( n5637 , n40 );
and ( n5638 , n5636 , n5637 );
not ( n5639 , n5222 );
or ( n5640 , n5639 , n5347 );
not ( n5641 , n5221 );
nor ( n5642 , n5352 , n5641 );
nand ( n5643 , n5640 , n5642 );
and ( n5644 , n844 , n5643 );
nor ( n5645 , n5638 , n5644 );
nand ( n5646 , n790 , n5186 );
nand ( n5647 , n5630 , n5645 , n5646 );
nor ( n5648 , n5625 , n5647 );
not ( n5649 , n5518 );
or ( n5650 , n5635 , n5649 );
not ( n5651 , n5362 );
and ( n5652 , n5651 , n5057 );
buf ( n5653 , n4937 );
and ( n5654 , n5359 , n5653 );
nor ( n5655 , n5652 , n5654 );
not ( n5656 , n4892 );
and ( n5657 , n5656 , n782 , n5361 );
nor ( n5658 , n5657 , n5371 );
nand ( n5659 , n5650 , n5655 , n5658 );
and ( n5660 , n40 , n5659 );
and ( n5661 , n848 , n5222 );
and ( n5662 , n5325 , n4429 );
not ( n5663 , n4686 );
and ( n5664 , n5322 , n5663 );
nor ( n5665 , n5662 , n5664 );
and ( n5666 , n5348 , n5624 );
nor ( n5667 , n5666 , n5332 );
nand ( n5668 , n5665 , n5667 );
and ( n5669 , n856 , n5668 );
nor ( n5670 , n5660 , n5661 , n5669 );
nand ( n5671 , n5648 , n5411 , n5670 );
nand ( n5672 , n2183 , n5671 );
and ( n5673 , n440 , n5624 );
not ( n5674 , n20 );
and ( n5675 , n5674 , n5431 );
nor ( n5676 , n5673 , n5675 , n5581 );
not ( n5677 , n288 );
and ( n5678 , n5677 , n5636 );
and ( n5679 , n2232 , n5643 );
nor ( n5680 , n5433 , n5430 );
and ( n5681 , n454 , n5680 );
nor ( n5682 , n5678 , n5679 , n5681 );
not ( n5683 , n2256 );
not ( n5684 , n5629 );
and ( n5685 , n5683 , n5684 );
and ( n5686 , n2268 , n5186 );
nor ( n5687 , n5685 , n5686 );
not ( n5688 , n40 );
and ( n5689 , n5688 , n5659 );
and ( n5690 , n445 , n5689 );
not ( n5691 , n2270 );
not ( n5692 , n5222 );
or ( n5693 , n5691 , n5692 );
not ( n5694 , n2199 );
nand ( n5695 , n5694 , n5668 );
nand ( n5696 , n5693 , n5695 );
nor ( n5697 , n5690 , n5696 );
nand ( n5698 , n5676 , n5682 , n5687 , n5697 );
nand ( n5699 , n2121 , n5698 );
not ( n5700 , n2 );
nand ( n5701 , n5700 , n5307 );
nand ( n5702 , n5617 , n5672 , n5699 , n5701 );
nor ( n5703 , n5606 , n5702 );
and ( n5704 , n2636 , n5636 );
not ( n5705 , n2681 );
nand ( n5706 , n5103 , n5705 );
not ( n5707 , n5328 );
and ( n5708 , n2308 , n5707 );
not ( n5709 , n2308 );
not ( n5710 , n23 );
and ( n5711 , n5709 , n5710 );
or ( n5712 , n5708 , n5711 );
or ( n5713 , n5706 , n5712 );
nor ( n5714 , n17 , n5712 );
nor ( n5715 , n15 , n5712 );
and ( n5716 , n2347 , n5715 );
or ( n5717 , n5714 , n5716 );
and ( n5718 , n2679 , n5717 );
and ( n5719 , n454 , n5716 );
nor ( n5720 , n5718 , n5719 );
nand ( n5721 , n5713 , n5720 );
not ( n5722 , n2664 );
not ( n5723 , n5643 );
or ( n5724 , n5722 , n5723 );
not ( n5725 , n2608 );
nand ( n5726 , n5725 , n5624 );
nand ( n5727 , n5724 , n5726 );
nor ( n5728 , n5704 , n5721 , n5727 );
not ( n5729 , n5712 );
and ( n5730 , n5729 , n2193 , n5103 );
not ( n5731 , n2675 );
not ( n5732 , n5186 );
or ( n5733 , n5731 , n5732 );
or ( n5734 , n2666 , n5629 );
nand ( n5735 , n5733 , n5734 );
nor ( n5736 , n5730 , n5735 );
and ( n5737 , n41 , n5689 );
not ( n5738 , n2671 );
not ( n5739 , n5668 );
or ( n5740 , n5738 , n5739 );
or ( n5741 , n2688 , n5639 );
nand ( n5742 , n5740 , n5741 );
nor ( n5743 , n5737 , n5742 );
and ( n5744 , n5728 , n5736 , n5743 );
nor ( n5745 , n5744 , n2662 );
not ( n5746 , n2697 );
not ( n5747 , n5239 );
or ( n5748 , n5746 , n5747 );
or ( n5749 , n2654 , n5441 );
and ( n5750 , n5487 , n41 );
and ( n5751 , n2630 , n5163 );
nor ( n5752 , n5750 , n5751 );
and ( n5753 , n2645 , n5460 );
and ( n5754 , n2633 , n5465 );
nor ( n5755 , n5753 , n5754 );
nand ( n5756 , n5749 , n5752 , n5755 );
not ( n5757 , n20 );
nand ( n5758 , n5729 , n5103 , n4074 );
or ( n5759 , n5757 , n5758 );
and ( n5760 , n5729 , n908 , n5103 );
not ( n5761 , n14 );
nor ( n5762 , n5712 , n5761 , n5405 );
and ( n5763 , n2066 , n5762 );
nor ( n5764 , n5760 , n5763 );
nand ( n5765 , n2719 , n5421 );
nand ( n5766 , n5759 , n5764 , n5765 );
or ( n5767 , n5756 , n5766 );
nand ( n5768 , n5767 , n2580 );
nand ( n5769 , n5748 , n5768 );
nor ( n5770 , n5745 , n5769 );
not ( n5771 , n2662 );
not ( n5772 , n5539 );
or ( n5773 , n5772 , n445 );
or ( n5774 , n2704 , n5549 );
nand ( n5775 , n5773 , n5774 );
not ( n5776 , n2630 );
not ( n5777 , n5217 );
or ( n5778 , n5776 , n5777 );
or ( n5779 , n2654 , n5522 );
nand ( n5780 , n5778 , n5779 );
nor ( n5781 , n5775 , n5780 );
or ( n5782 , n2637 , n5516 );
nand ( n5783 , n5781 , n5764 , n5782 , n5759 );
nand ( n5784 , n5771 , n5783 );
not ( n5785 , n2604 );
not ( n5786 , n5758 );
and ( n5787 , n5785 , n5786 );
nor ( n5788 , n5712 , n5405 , n2596 );
nor ( n5789 , n5787 , n5788 );
and ( n5790 , n2609 , n5320 );
not ( n5791 , n2592 );
and ( n5792 , n5791 , n5762 );
nor ( n5793 , n5790 , n5792 );
and ( n5794 , n5770 , n5784 , n5789 , n5793 );
and ( n5795 , n5495 , n5703 , n5794 );
nand ( n5796 , n1 , n4254 );
nor ( n5797 , n5795 , n5796 );
not ( n5798 , n3371 );
not ( n5799 , n3516 );
nor ( n5800 , n5799 , n5409 );
and ( n5801 , n3609 , n5798 , n5800 );
not ( n5802 , n4380 );
nand ( n5803 , n5802 , n5048 );
or ( n5804 , n3371 , n3874 , n5803 );
not ( n5805 , n40 );
or ( n5806 , n5805 , n31 );
not ( n5807 , n3604 );
or ( n5808 , n40 , n5807 );
nand ( n5809 , n5806 , n5808 , n23 );
or ( n5810 , n4214 , n5809 );
nand ( n5811 , n5804 , n5810 );
nor ( n5812 , n5801 , n5811 );
not ( n5813 , n13 );
nand ( n5814 , n5813 , n3516 );
not ( n5815 , n5814 );
not ( n5816 , n3813 );
not ( n5817 , n5816 );
not ( n5818 , n5817 );
not ( n5819 , n5818 );
not ( n5820 , n5819 );
not ( n5821 , n5820 );
not ( n5822 , n5821 );
nor ( n5823 , n3609 , n5822 );
nand ( n5824 , n5815 , n5823 , n3119 , n2056 );
not ( n5825 , n5814 );
nand ( n5826 , n23 , n3575 );
not ( n5827 , n5826 );
not ( n5828 , n5827 );
not ( n5829 , n5828 );
not ( n5830 , n5829 );
nor ( n5831 , n3609 , n5830 );
not ( n5832 , n290 );
nand ( n5833 , n5825 , n3119 , n5831 , n5832 );
not ( n5834 , n13 );
not ( n5835 , n3516 );
nand ( n5836 , n5834 , n5835 );
not ( n5837 , n5830 );
not ( n5838 , n5837 );
nand ( n5839 , n5838 , n5803 );
and ( n5840 , n287 , n5839 );
nand ( n5841 , n5822 , n5803 );
and ( n5842 , n286 , n5841 );
nor ( n5843 , n5840 , n5842 );
nor ( n5844 , n5836 , n5843 );
nand ( n5845 , n39 , n985 , n5844 );
and ( n5846 , n5812 , n5824 , n5833 , n5845 );
not ( n5847 , n2781 );
not ( n5848 , n23 );
nand ( n5849 , n5848 , n5803 );
not ( n5850 , n5849 );
not ( n5851 , n5850 );
nand ( n5852 , n5847 , n5851 );
or ( n5853 , n39 , n5852 );
not ( n5854 , n5839 );
or ( n5855 , n3874 , n5854 );
and ( n5856 , n2781 , n5831 );
and ( n5857 , n3609 , n5149 );
nor ( n5858 , n5856 , n5857 );
nand ( n5859 , n5853 , n5855 , n5858 );
and ( n5860 , n994 , n5859 );
not ( n5861 , n3368 );
nor ( n5862 , n3493 , n5861 );
not ( n5863 , n5862 );
nand ( n5864 , n5329 , n5803 );
and ( n5865 , n40 , n5864 );
not ( n5866 , n40 );
and ( n5867 , n5866 , n5849 );
nor ( n5868 , n5865 , n5867 );
nor ( n5869 , n5863 , n5868 );
and ( n5870 , n3609 , n5869 );
nor ( n5871 , n5860 , n5870 );
nand ( n5872 , n3609 , n985 );
not ( n5873 , n5571 );
nor ( n5874 , n5873 , n5575 );
or ( n5875 , n13 , n5872 , n5874 );
not ( n5876 , n2579 );
not ( n5877 , n5858 );
and ( n5878 , n5876 , n5877 );
and ( n5879 , n1849 , n5859 );
nor ( n5880 , n5878 , n5879 );
nand ( n5881 , n2898 , n5049 );
not ( n5882 , n5881 );
buf ( n5883 , n5882 );
not ( n5884 , n5883 );
buf ( n5885 , n5884 );
not ( n5886 , n5885 );
nor ( n5887 , n2616 , n5886 );
and ( n5888 , n5887 , n5282 );
not ( n5889 , n5837 );
nor ( n5890 , n5889 , n1995 );
not ( n5891 , n5890 );
not ( n5892 , n5883 );
and ( n5893 , n1938 , n5892 );
nand ( n5894 , n5167 , n5893 , n5292 );
nand ( n5895 , n5891 , n5894 );
nor ( n5896 , n5888 , n5895 );
nand ( n5897 , n23 , n5826 );
not ( n5898 , n5897 );
not ( n5899 , n5898 );
not ( n5900 , n5899 );
not ( n5901 , n5900 );
not ( n5902 , n5901 );
not ( n5903 , n5902 );
not ( n5904 , n5903 );
not ( n5905 , n5882 );
and ( n5906 , n5167 , n5905 , n4390 );
not ( n5907 , n23 );
not ( n5908 , n24 );
nor ( n5909 , n5908 , n22 );
nand ( n5910 , n5909 , n5063 , n5048 );
nand ( n5911 , n5907 , n5910 );
nor ( n5912 , n5906 , n5911 );
or ( n5913 , n5166 , n5912 );
not ( n5914 , n5253 );
and ( n5915 , n5171 , n5905 , n5914 );
nor ( n5916 , n5915 , n5911 );
or ( n5917 , n795 , n5916 );
nand ( n5918 , n5913 , n5917 );
not ( n5919 , n5918 );
or ( n5920 , n5904 , n5919 );
nor ( n5921 , n19 , n5889 );
nand ( n5922 , n724 , n5921 );
nand ( n5923 , n5920 , n5922 );
not ( n5924 , n5902 );
nand ( n5925 , n5924 , n2615 );
not ( n5926 , n5881 );
not ( n5927 , n5926 );
buf ( n5928 , n5927 );
not ( n5929 , n5928 );
or ( n5930 , n5929 , n4746 );
not ( n5931 , n5911 );
nand ( n5932 , n5930 , n5931 );
not ( n5933 , n5932 );
or ( n5934 , n5925 , n5933 );
not ( n5935 , n5927 );
nor ( n5936 , n795 , n5935 );
nand ( n5937 , n5171 , n5936 , n5254 );
nand ( n5938 , n5934 , n5937 );
nor ( n5939 , n5923 , n5938 );
nand ( n5940 , n5896 , n5939 );
and ( n5941 , n5940 , n3629 , n1982 );
or ( n5942 , n2616 , n5933 );
nand ( n5943 , n5942 , n5919 );
and ( n5944 , n3609 , n3069 , n5943 );
nor ( n5945 , n5941 , n5944 );
nand ( n5946 , n5880 , n5945 );
nand ( n5947 , n3609 , n1982 );
not ( n5948 , n914 );
not ( n5949 , n5884 );
or ( n5950 , n5949 , n5152 );
nand ( n5951 , n5950 , n5931 );
not ( n5952 , n5951 );
or ( n5953 , n5948 , n5952 );
or ( n5954 , n5093 , n5935 , n4995 );
nand ( n5955 , n5954 , n5931 );
and ( n5956 , n909 , n5955 );
not ( n5957 , n5881 );
nor ( n5958 , n4318 , n5957 );
or ( n5959 , n5911 , n5958 );
and ( n5960 , n942 , n5959 );
nor ( n5961 , n5956 , n5960 );
nand ( n5962 , n5953 , n5961 );
or ( n5963 , n5929 , n4933 );
nand ( n5964 , n5963 , n5931 );
not ( n5965 , n5964 );
or ( n5966 , n765 , n5965 );
or ( n5967 , n5949 , n4872 );
nand ( n5968 , n5967 , n5931 );
not ( n5969 , n5968 );
or ( n5970 , n585 , n5969 );
not ( n5971 , n782 );
and ( n5972 , n5927 , n5109 );
nor ( n5973 , n5972 , n5911 );
or ( n5974 , n5971 , n5973 );
nand ( n5975 , n5966 , n5970 , n5974 );
nor ( n5976 , n5962 , n5975 );
or ( n5977 , n5947 , n5976 );
or ( n5978 , n3664 , n3501 );
not ( n5979 , n5903 );
not ( n5980 , n5979 );
not ( n5981 , n5980 );
not ( n5982 , n5981 );
nand ( n5983 , n5885 , n5082 );
nand ( n5984 , n5931 , n5983 );
and ( n5985 , n5982 , n5984 );
not ( n5986 , n5838 );
not ( n5987 , n5986 );
nand ( n5988 , n5987 , n5983 );
nor ( n5989 , n5985 , n5988 );
or ( n5990 , n5978 , n5989 );
not ( n5991 , n5243 );
nor ( n5992 , n5886 , n5991 );
and ( n5993 , n97 , n5992 );
not ( n5994 , n5890 );
nand ( n5995 , n4423 , n5893 , n5257 );
nand ( n5996 , n5994 , n5995 );
not ( n5997 , n5288 );
and ( n5998 , n5285 , n5936 , n5997 );
nor ( n5999 , n5993 , n5996 , n5998 );
not ( n6000 , n97 );
not ( n6001 , n5928 );
or ( n6002 , n6001 , n5242 );
nand ( n6003 , n6002 , n5931 );
not ( n6004 , n6003 );
or ( n6005 , n6000 , n6004 );
not ( n6006 , n4423 );
or ( n6007 , n6006 , n5883 , n4417 );
nand ( n6008 , n6007 , n5931 );
and ( n6009 , n2125 , n6008 );
or ( n6010 , n5284 , n5883 , n5286 );
nand ( n6011 , n6010 , n5931 );
and ( n6012 , n2123 , n6011 );
nor ( n6013 , n6009 , n6012 );
nand ( n6014 , n6005 , n6013 );
and ( n6015 , n5980 , n6014 );
and ( n6016 , n96 , n5921 );
nor ( n6017 , n6015 , n6016 );
nand ( n6018 , n5999 , n6017 );
nand ( n6019 , n2603 , n6018 );
or ( n6020 , n3609 , n6019 );
nand ( n6021 , n5977 , n5990 , n6020 );
nor ( n6022 , n5946 , n6021 );
nand ( n6023 , n39 , n1982 );
not ( n6024 , n6023 );
not ( n6025 , n5979 );
and ( n6026 , n5962 , n6025 );
not ( n6027 , n5928 );
nor ( n6028 , n913 , n6027 );
and ( n6029 , n6028 , n5482 );
nor ( n6030 , n5828 , n521 );
and ( n6031 , n908 , n6030 );
nor ( n6032 , n6026 , n6029 , n6031 );
nor ( n6033 , n912 , n5838 , n633 );
not ( n6034 , n6033 );
not ( n6035 , n6027 );
nand ( n6036 , n909 , n6035 );
nor ( n6037 , n6036 , n4995 );
and ( n6038 , n6037 , n5028 );
and ( n6039 , n942 , n5958 );
nor ( n6040 , n6038 , n6039 );
nand ( n6041 , n6032 , n6034 , n6040 );
and ( n6042 , n6024 , n6041 );
not ( n6043 , n5984 );
nor ( n6044 , n3501 , n6043 );
and ( n6045 , n3664 , n6044 );
and ( n6046 , n5980 , n5975 );
nor ( n6047 , n765 , n5886 );
not ( n6048 , n6047 );
not ( n6049 , n5262 );
or ( n6050 , n6048 , n6049 );
nor ( n6051 , n585 , n6027 );
not ( n6052 , n5265 );
and ( n6053 , n6051 , n6052 );
or ( n6054 , n6027 , n5365 );
and ( n6055 , n2457 , n5829 , n5368 );
and ( n6056 , n624 , n6030 );
nor ( n6057 , n6055 , n6056 );
nand ( n6058 , n6054 , n6057 );
nor ( n6059 , n6053 , n6058 );
nand ( n6060 , n6050 , n6059 );
nor ( n6061 , n6046 , n6060 );
or ( n6062 , n6023 , n6061 );
nand ( n6063 , n5928 , n5161 );
nand ( n6064 , n5931 , n6063 );
nand ( n6065 , n6064 , n3069 , n3643 );
nand ( n6066 , n6062 , n6065 );
nor ( n6067 , n6042 , n6045 , n6066 );
not ( n6068 , n6014 );
not ( n6069 , n6068 );
and ( n6070 , n3609 , n2603 , n6069 );
and ( n6071 , n5980 , n6064 );
not ( n6072 , n5986 );
nand ( n6073 , n6072 , n6063 );
nor ( n6074 , n6071 , n6073 );
nor ( n6075 , n6074 , n3070 , n3645 );
nor ( n6076 , n6070 , n6075 );
not ( n6077 , n6035 );
not ( n6078 , n4937 );
or ( n6079 , n6077 , n6078 );
nand ( n6080 , n6079 , n5931 );
not ( n6081 , n6080 );
or ( n6082 , n765 , n6081 );
or ( n6083 , n5886 , n4876 );
nand ( n6084 , n6083 , n5931 );
and ( n6085 , n584 , n6084 );
nor ( n6086 , n5926 , n4892 );
nor ( n6087 , n6086 , n5911 );
nor ( n6088 , n6087 , n5971 );
nor ( n6089 , n6085 , n6088 );
nand ( n6090 , n6082 , n6089 );
and ( n6091 , n3609 , n6090 );
not ( n6092 , n20 );
not ( n6093 , n3664 );
not ( n6094 , n6027 );
nand ( n6095 , n6094 , n4585 );
nand ( n6096 , n5931 , n6095 );
not ( n6097 , n6096 );
or ( n6098 , n6093 , n6097 );
nand ( n6099 , n6098 , n5858 );
and ( n6100 , n6092 , n6099 );
nor ( n6101 , n6091 , n6100 );
not ( n6102 , n2615 );
not ( n6103 , n6096 );
not ( n6104 , n5980 );
or ( n6105 , n6103 , n6104 );
not ( n6106 , n5986 );
and ( n6107 , n6106 , n6095 );
nand ( n6108 , n6105 , n6107 );
not ( n6109 , n6108 );
or ( n6110 , n6102 , n6109 );
not ( n6111 , n4428 );
and ( n6112 , n5893 , n6111 );
and ( n6113 , n5936 , n5663 );
nor ( n6114 , n6112 , n6113 );
not ( n6115 , n14 );
and ( n6116 , n5663 , n5905 );
nor ( n6117 , n6116 , n5911 );
and ( n6118 , n6115 , n6117 );
and ( n6119 , n5927 , n4427 );
nor ( n6120 , n6119 , n5911 );
and ( n6121 , n14 , n6120 );
nor ( n6122 , n6118 , n6121 , n432 );
and ( n6123 , n6025 , n6122 );
nor ( n6124 , n6123 , n5890 );
and ( n6125 , n6114 , n6124 );
nand ( n6126 , n6110 , n6125 );
and ( n6127 , n3659 , n6126 );
nand ( n6128 , n6035 , n4816 );
nand ( n6129 , n5931 , n6128 );
nand ( n6130 , n5980 , n6129 );
not ( n6131 , n6128 );
nor ( n6132 , n5986 , n6131 );
nand ( n6133 , n6130 , n6132 );
and ( n6134 , n3646 , n6133 );
nor ( n6135 , n6127 , n6134 );
and ( n6136 , n97 , n6129 );
nor ( n6137 , n6136 , n6122 );
not ( n6138 , n6137 );
nand ( n6139 , n6138 , n3735 );
not ( n6140 , n5981 );
not ( n6141 , n1571 );
not ( n6142 , n6080 );
or ( n6143 , n6141 , n6142 );
nand ( n6144 , n6143 , n6089 );
and ( n6145 , n6140 , n6144 );
and ( n6146 , n6047 , n5653 );
nor ( n6147 , n6145 , n6146 );
nand ( n6148 , n782 , n6086 );
and ( n6149 , n6051 , n5057 );
not ( n6150 , n6057 );
nor ( n6151 , n6149 , n6150 );
nand ( n6152 , n6147 , n6148 , n6151 );
nand ( n6153 , n39 , n6152 );
nand ( n6154 , n6101 , n6135 , n6139 , n6153 );
and ( n6155 , n2517 , n6154 );
not ( n6156 , n3643 );
nand ( n6157 , n6094 , n4670 );
nand ( n6158 , n5931 , n6157 );
not ( n6159 , n6158 );
or ( n6160 , n6156 , n6159 );
nand ( n6161 , n5980 , n6158 );
and ( n6162 , n6161 , n5987 , n6157 );
or ( n6163 , n6162 , n3645 );
nand ( n6164 , n6160 , n6163 );
and ( n6165 , n20 , n6164 );
not ( n6166 , n3629 );
not ( n6167 , n6094 );
not ( n6168 , n4750 );
or ( n6169 , n6167 , n6168 );
nand ( n6170 , n6169 , n5931 );
not ( n6171 , n6170 );
or ( n6172 , n6171 , n5925 );
nand ( n6173 , n6172 , n5922 );
not ( n6174 , n6173 );
and ( n6175 , n5887 , n4750 );
nor ( n6176 , n6175 , n5890 );
nand ( n6177 , n5936 , n4480 );
not ( n6178 , n5904 );
or ( n6179 , n5926 , n4397 );
nand ( n6180 , n6179 , n5931 );
and ( n6181 , n14 , n6180 );
not ( n6182 , n14 );
or ( n6183 , n5926 , n4479 );
nand ( n6184 , n6183 , n5931 );
and ( n6185 , n6182 , n6184 );
nor ( n6186 , n6181 , n6185 );
nor ( n6187 , n6186 , n432 );
and ( n6188 , n6178 , n6187 );
and ( n6189 , n5893 , n4398 );
nor ( n6190 , n6188 , n6189 );
nand ( n6191 , n6174 , n6176 , n6177 , n6190 );
not ( n6192 , n6191 );
or ( n6193 , n6166 , n6192 );
not ( n6194 , n2615 );
not ( n6195 , n6170 );
or ( n6196 , n6194 , n6195 );
not ( n6197 , n6187 );
nand ( n6198 , n6196 , n6197 );
nand ( n6199 , n20 , n6198 );
not ( n6200 , n6199 );
nand ( n6201 , n3609 , n6200 );
nand ( n6202 , n6193 , n6201 );
nor ( n6203 , n6165 , n6202 );
and ( n6204 , n6028 , n4990 );
nor ( n6205 , n6204 , n6033 );
not ( n6206 , n5987 );
nand ( n6207 , n6206 , n909 );
not ( n6208 , n5931 );
nand ( n6209 , n5885 , n4326 );
not ( n6210 , n6209 );
or ( n6211 , n6208 , n6210 );
nand ( n6212 , n6211 , n942 );
or ( n6213 , n6027 , n4989 );
nand ( n6214 , n6213 , n5931 );
and ( n6215 , n914 , n6214 );
nand ( n6216 , n5885 , n5029 );
and ( n6217 , n5931 , n6216 );
nor ( n6218 , n6217 , n910 );
nor ( n6219 , n6215 , n6218 );
nand ( n6220 , n6212 , n6219 );
and ( n6221 , n6140 , n6220 );
or ( n6222 , n6036 , n5030 );
or ( n6223 , n963 , n6209 );
nand ( n6224 , n6222 , n6223 );
nor ( n6225 , n6221 , n6224 );
nand ( n6226 , n6205 , n6207 , n6225 );
and ( n6227 , n39 , n6226 );
not ( n6228 , n6220 );
or ( n6229 , n39 , n6228 );
not ( n6230 , n20 );
or ( n6231 , n6230 , n5858 );
nand ( n6232 , n6229 , n6231 );
nor ( n6233 , n6227 , n6232 );
and ( n6234 , n6203 , n6233 );
not ( n6235 , n2517 );
nor ( n6236 , n6234 , n6235 );
nor ( n6237 , n6155 , n6236 );
nand ( n6238 , n6022 , n6067 , n6076 , n6237 );
not ( n6239 , n2 );
and ( n6240 , n6238 , n6239 );
and ( n6241 , n87 , n5864 );
not ( n6242 , n87 );
and ( n6243 , n6242 , n5849 );
nor ( n6244 , n6241 , n6243 );
not ( n6245 , n6244 );
not ( n6246 , n6245 );
nor ( n6247 , n6246 , n5836 , n5872 );
nor ( n6248 , n6240 , n6247 );
and ( n6249 , n5846 , n5871 , n5875 , n6248 );
or ( n6250 , n6249 , n3751 );
nand ( n6251 , n4 , n5 );
nand ( n6252 , n3 , n3569 );
nand ( n6253 , n6251 , n6252 );
not ( n6254 , n6253 );
not ( n6255 , n2 );
not ( n6256 , n908 );
nor ( n6257 , n5033 , n5405 );
not ( n6258 , n6257 );
or ( n6259 , n6256 , n6258 );
nand ( n6260 , n6259 , n6228 );
and ( n6261 , n2517 , n6260 );
not ( n6262 , n5951 );
or ( n6263 , n632 , n6262 );
and ( n6264 , n520 , n5955 );
nor ( n6265 , n6264 , n6257 );
nand ( n6266 , n6263 , n6265 );
and ( n6267 , n2041 , n6266 );
nor ( n6268 , n6261 , n6267 );
nand ( n6269 , n4881 , n5103 );
nand ( n6270 , n583 , n5968 );
and ( n6271 , n6269 , n6270 );
and ( n6272 , n764 , n5964 );
nor ( n6273 , n1375 , n5973 );
nor ( n6274 , n6272 , n6273 );
nand ( n6275 , n6271 , n6274 );
nand ( n6276 , n6275 , n1984 , n1982 );
not ( n6277 , n2617 );
not ( n6278 , n6096 );
or ( n6279 , n6277 , n6278 );
nand ( n6280 , n453 , n5149 );
nand ( n6281 , n6279 , n6280 );
or ( n6282 , n3264 , n6120 );
or ( n6283 , n20 , n795 );
or ( n6284 , n6283 , n6117 );
not ( n6285 , n20 );
nand ( n6286 , n6285 , n97 );
not ( n6287 , n6286 );
nand ( n6288 , n6287 , n6129 );
not ( n6289 , n20 );
and ( n6290 , n764 , n6080 );
nor ( n6291 , n6087 , n1375 );
nor ( n6292 , n6290 , n6291 );
nand ( n6293 , n583 , n6084 );
nand ( n6294 , n6292 , n6269 , n6293 );
nand ( n6295 , n6289 , n6294 );
nand ( n6296 , n6282 , n6284 , n6288 , n6295 );
or ( n6297 , n6281 , n6296 );
nand ( n6298 , n6297 , n2517 );
and ( n6299 , n6268 , n6276 , n6298 );
or ( n6300 , n3425 , n1314 );
nand ( n6301 , n6300 , n4330 );
or ( n6302 , n6301 , n5405 , n1971 );
or ( n6303 , n2579 , n6280 );
nand ( n6304 , n6302 , n6303 );
or ( n6305 , n3454 , n1971 , n5104 );
not ( n6306 , n5959 );
or ( n6307 , n1990 , n6306 );
nand ( n6308 , n6305 , n6307 );
nor ( n6309 , n6304 , n6308 );
or ( n6310 , n1316 , n6171 );
not ( n6311 , n6158 );
or ( n6312 , n295 , n6311 );
nand ( n6313 , n6310 , n6312 );
and ( n6314 , n6313 , n1852 , n1314 );
nand ( n6315 , n5104 , n5852 );
and ( n6316 , n1849 , n6315 );
nor ( n6317 , n6314 , n6316 );
and ( n6318 , n2018 , n6008 );
and ( n6319 , n1998 , n6011 );
nor ( n6320 , n6318 , n6319 );
and ( n6321 , n1985 , n5918 );
nor ( n6322 , n6197 , n3471 , n1971 );
nor ( n6323 , n6321 , n6322 );
and ( n6324 , n2030 , n6064 );
nor ( n6325 , n6324 , n6044 );
and ( n6326 , n3482 , n6003 );
and ( n6327 , n2014 , n5932 );
nor ( n6328 , n6326 , n6327 );
and ( n6329 , n6320 , n6323 , n6325 , n6328 );
nand ( n6330 , n6299 , n6309 , n6317 , n6329 );
and ( n6331 , n6255 , n6330 );
nor ( n6332 , n6246 , n3516 , n81 );
nor ( n6333 , n6331 , n6332 );
not ( n6334 , n5864 );
and ( n6335 , n2310 , n6334 );
not ( n6336 , n2310 );
and ( n6337 , n6336 , n5850 );
or ( n6338 , n6335 , n6337 );
not ( n6339 , n6338 );
not ( n6340 , n3516 );
and ( n6341 , n6339 , n6340 , n3531 );
nor ( n6342 , n6341 , n5869 );
and ( n6343 , n3525 , n6315 );
not ( n6344 , n3531 );
nor ( n6345 , n5405 , n6344 );
and ( n6346 , n6345 , n5729 );
or ( n6347 , n81 , n5430 );
or ( n6348 , n5409 , n3369 );
nand ( n6349 , n6347 , n6348 );
and ( n6350 , n5103 , n6349 );
nor ( n6351 , n6343 , n6346 , n6350 );
nand ( n6352 , n6333 , n6342 , n6351 );
not ( n6353 , n6352 );
or ( n6354 , n6254 , n6353 );
not ( n6355 , n4253 );
or ( n6356 , n6338 , n42 );
nand ( n6357 , n42 , n5729 );
nand ( n6358 , n6356 , n6357 );
and ( n6359 , n942 , n6358 );
not ( n6360 , n2389 );
or ( n6361 , n2396 , n6338 );
and ( n6362 , n2398 , n5729 );
and ( n6363 , n17 , n5715 );
nor ( n6364 , n6362 , n6363 );
nand ( n6365 , n6361 , n6364 );
not ( n6366 , n6365 );
nor ( n6367 , n6360 , n6366 );
or ( n6368 , n2387 , n2384 );
nand ( n6369 , n6368 , n2391 );
nand ( n6370 , n6369 , n6365 );
not ( n6371 , n6370 );
nor ( n6372 , n2493 , n5279 );
or ( n6373 , n6359 , n6367 , n6371 , n6372 );
not ( n6374 , n6373 );
and ( n6375 , n5285 , n2418 , n5289 );
nor ( n6376 , n5248 , n841 , n2501 );
nor ( n6377 , n6375 , n6376 );
nand ( n6378 , n2463 , n4890 );
not ( n6379 , n6378 );
nand ( n6380 , n5729 , n5103 , n1919 );
and ( n6381 , n5171 , n2802 , n5254 );
nand ( n6382 , n20 , n6381 );
nand ( n6383 , n2409 , n4319 );
or ( n6384 , n2306 , n6338 );
and ( n6385 , n2332 , n5717 );
not ( n6386 , n6357 );
and ( n6387 , n2123 , n6386 );
nor ( n6388 , n6385 , n6387 );
nand ( n6389 , n6384 , n6388 );
nand ( n6390 , n20 , n6389 );
nand ( n6391 , n6380 , n6382 , n6383 , n6390 );
nor ( n6392 , n4378 , n2431 , n5293 );
nor ( n6393 , n6006 , n3182 , n5258 );
nor ( n6394 , n6379 , n6391 , n6392 , n6393 );
or ( n6395 , n912 , n2498 , n4995 , n5093 );
nand ( n6396 , n6374 , n6377 , n6394 , n6395 );
and ( n6397 , n724 , n6358 );
and ( n6398 , n16 , n5717 );
nor ( n6399 , n6397 , n6398 );
nor ( n6400 , n2435 , n6399 );
and ( n6401 , n520 , n6358 );
not ( n6402 , n16 );
and ( n6403 , n6402 , n5717 );
nor ( n6404 , n6401 , n6403 );
nor ( n6405 , n912 , n6404 );
nor ( n6406 , n6396 , n6400 , n6405 );
and ( n6407 , n2468 , n6365 );
or ( n6408 , n841 , n6399 );
or ( n6409 , n2242 , n6366 );
and ( n6410 , n5729 , n5103 , n3345 );
and ( n6411 , n570 , n6358 );
nor ( n6412 , n6410 , n6411 );
nand ( n6413 , n6408 , n6409 , n6412 );
not ( n6414 , n2478 );
nor ( n6415 , n6414 , n5244 );
not ( n6416 , n6415 );
not ( n6417 , n20 );
nand ( n6418 , n6417 , n6389 );
not ( n6419 , n6052 );
not ( n6420 , n6419 );
nand ( n6421 , n3350 , n6420 );
or ( n6422 , n3176 , n6404 );
nand ( n6423 , n6416 , n6418 , n6421 , n6422 );
nor ( n6424 , n6407 , n6413 , n6423 );
nand ( n6425 , n2475 , n5262 );
not ( n6426 , n6368 );
and ( n6427 , n5482 , n2398 , n6426 );
nor ( n6428 , n4746 , n645 , n2501 );
nor ( n6429 , n6427 , n6428 );
nand ( n6430 , n6406 , n6424 , n6425 , n6429 );
nand ( n6431 , n6355 , n1982 , n2508 , n6430 );
nand ( n6432 , n6354 , n6431 );
not ( n6433 , n6432 );
nand ( n6434 , n4194 , n5859 );
nand ( n6435 , n6250 , n6433 , n6434 );
nor ( n6436 , n5797 , n6435 );
nor ( n6437 , n3118 , n2731 );
and ( n6438 , n5844 , n3937 , n6437 );
not ( n6439 , n2299 );
and ( n6440 , n4158 , n1852 );
not ( n6441 , n6440 );
nor ( n6442 , n5715 , n5714 );
nor ( n6443 , n6439 , n6441 , n6442 , n38 );
nor ( n6444 , n6438 , n6443 );
nand ( n6445 , n1980 , n3798 );
or ( n6446 , n13 , n6445 , n2731 , n5874 );
and ( n6447 , n4184 , n5862 );
nand ( n6448 , n3609 , n5839 );
or ( n6449 , n40 , n6448 );
or ( n6450 , n3609 , n5868 );
nand ( n6451 , n40 , n3609 );
not ( n6452 , n5841 );
or ( n6453 , n6451 , n6452 );
nand ( n6454 , n6449 , n6450 , n6453 );
nand ( n6455 , n38 , n2298 , n6447 , n6454 );
and ( n6456 , n6444 , n6446 , n6455 );
not ( n6457 , n3516 );
nand ( n6458 , n2299 , n6457 );
nor ( n6459 , n6458 , n6338 );
and ( n6460 , n6459 , n3938 , n6440 );
not ( n6461 , n6440 );
and ( n6462 , n2576 , n5839 );
and ( n6463 , n2577 , n5841 );
nor ( n6464 , n6462 , n6463 );
nor ( n6465 , n6461 , n6458 , n6464 , n3938 );
nor ( n6466 , n6460 , n6465 );
not ( n6467 , n2889 );
not ( n6468 , n6352 );
or ( n6469 , n6467 , n6468 );
or ( n6470 , n3766 , n5852 );
and ( n6471 , n3771 , n5839 );
not ( n6472 , n17 );
nor ( n6473 , n15 , n39 );
and ( n6474 , n38 , n6473 , n5827 );
not ( n6475 , n23 );
nor ( n6476 , n6475 , n15 );
and ( n6477 , n3763 , n6476 );
nor ( n6478 , n6474 , n6477 );
or ( n6479 , n6472 , n6478 );
and ( n6480 , n38 , n3882 , n5827 );
not ( n6481 , n23 );
nor ( n6482 , n6481 , n17 );
and ( n6483 , n3763 , n6482 );
nor ( n6484 , n6480 , n6483 );
nand ( n6485 , n6479 , n6484 );
nor ( n6486 , n6471 , n6485 );
nand ( n6487 , n6470 , n6486 );
nand ( n6488 , n6487 , n994 , n2301 );
nand ( n6489 , n6469 , n6488 );
not ( n6490 , n6489 );
nand ( n6491 , n6456 , n6466 , n6490 );
nor ( n6492 , n2 , n3 );
nand ( n6493 , n454 , n1982 );
not ( n6494 , n6493 );
or ( n6495 , n3789 , n6478 );
or ( n6496 , n14 , n6484 );
nand ( n6497 , n6495 , n6496 );
and ( n6498 , n6494 , n6497 );
or ( n6499 , n2244 , n6478 );
not ( n6500 , n14 );
or ( n6501 , n6500 , n6484 );
nand ( n6502 , n6499 , n6501 );
and ( n6503 , n3080 , n6502 );
nor ( n6504 , n6498 , n6503 );
and ( n6505 , n1849 , n6487 );
not ( n6506 , n2435 );
nand ( n6507 , n2234 , n6506 );
or ( n6508 , n6507 , n2579 );
nor ( n6509 , n2681 , n2579 );
not ( n6510 , n6509 );
nand ( n6511 , n6508 , n6510 );
and ( n6512 , n6511 , n6485 );
nor ( n6513 , n6505 , n6512 );
not ( n6514 , n3958 );
and ( n6515 , n5940 , n6514 , n1982 );
and ( n6516 , n5943 , n3934 , n3069 );
nor ( n6517 , n6515 , n6516 );
nor ( n6518 , n20 , n5947 );
and ( n6519 , n38 , n6518 , n6018 );
not ( n6520 , n6494 );
nor ( n6521 , n6520 , n2065 , n5989 , n3934 );
nor ( n6522 , n6519 , n6521 );
and ( n6523 , n6504 , n6513 , n6517 , n6522 );
nand ( n6524 , n3768 , n1982 );
or ( n6525 , n6524 , n6061 );
nand ( n6526 , n3769 , n3080 , n2229 , n6064 );
nand ( n6527 , n6525 , n6526 );
not ( n6528 , n3074 );
nor ( n6529 , n630 , n2579 );
not ( n6530 , n6529 );
and ( n6531 , n6528 , n6530 );
not ( n6532 , n6485 );
nor ( n6533 , n6531 , n6532 );
not ( n6534 , n3935 );
and ( n6535 , n6534 , n6494 , n450 , n5984 );
nor ( n6536 , n6527 , n6533 , n6535 );
not ( n6537 , n6524 );
and ( n6538 , n6537 , n6041 );
nor ( n6539 , n2579 , n3954 , n5976 );
nor ( n6540 , n6538 , n6539 );
nor ( n6541 , n2228 , n6074 );
and ( n6542 , n6541 , n3919 , n3080 );
and ( n6543 , n6069 , n3769 , n2603 );
nor ( n6544 , n6542 , n6543 );
and ( n6545 , n908 , n6485 );
and ( n6546 , n2066 , n6502 );
or ( n6547 , n6311 , n3766 , n2629 );
or ( n6548 , n6507 , n6532 );
nand ( n6549 , n6547 , n6548 );
nor ( n6550 , n6545 , n6546 , n6549 );
or ( n6551 , n2629 , n6162 );
not ( n6552 , n6226 );
nand ( n6553 , n6551 , n6552 );
and ( n6554 , n3919 , n6553 );
nand ( n6555 , n6199 , n6228 );
not ( n6556 , n6555 );
or ( n6557 , n3768 , n6556 );
not ( n6558 , n6191 );
or ( n6559 , n6558 , n3958 );
nand ( n6560 , n6557 , n6559 );
nor ( n6561 , n6554 , n6560 );
nand ( n6562 , n6550 , n6561 );
nand ( n6563 , n6562 , n2517 );
and ( n6564 , n454 , n6497 );
and ( n6565 , n2191 , n6485 );
nor ( n6566 , n6564 , n6565 );
and ( n6567 , n3943 , n6096 );
and ( n6568 , n5705 , n6485 );
nor ( n6569 , n6567 , n6568 );
and ( n6570 , n6566 , n6569 );
not ( n6571 , n3766 );
and ( n6572 , n6571 , n6144 );
not ( n6573 , n6108 );
or ( n6574 , n6573 , n3850 );
or ( n6575 , n3927 , n6125 );
nand ( n6576 , n6574 , n6575 );
nor ( n6577 , n6572 , n6576 );
not ( n6578 , n20 );
nand ( n6579 , n6578 , n3968 , n6133 );
not ( n6580 , n3842 );
not ( n6581 , n6137 );
and ( n6582 , n6580 , n6581 );
and ( n6583 , n3768 , n6152 );
nor ( n6584 , n6582 , n6583 );
nand ( n6585 , n6570 , n6577 , n6579 , n6584 );
nand ( n6586 , n2517 , n6585 );
and ( n6587 , n6544 , n6563 , n6586 );
nand ( n6588 , n6523 , n6536 , n6540 , n6587 );
nand ( n6589 , n6492 , n4184 , n6588 );
nand ( n6590 , n2299 , n3 , n6352 );
not ( n6591 , n4193 );
nand ( n6592 , n6591 , n2298 , n4184 );
not ( n6593 , n2 );
not ( n6594 , n6487 );
or ( n6595 , n6592 , n6593 , n6594 );
nand ( n6596 , n3920 , n6437 );
or ( n6597 , n6596 , n5836 , n6246 );
nand ( n6598 , n6595 , n6597 );
not ( n6599 , n6447 );
nor ( n6600 , n6599 , n3 , n38 , n5868 );
nand ( n6601 , n3936 , n2301 , n5798 , n5800 );
not ( n6602 , n5809 );
nand ( n6603 , n38 , n3516 );
nor ( n6604 , n39 , n6603 , n3371 );
nand ( n6605 , n6602 , n6604 , n2301 );
and ( n6606 , n39 , n5729 );
or ( n6607 , n3819 , n2575 );
nand ( n6608 , n6607 , n5822 );
and ( n6609 , n3609 , n6608 );
nor ( n6610 , n6606 , n6609 );
or ( n6611 , n6603 , n6441 , n5 , n6610 );
nor ( n6612 , n12 , n3832 );
not ( n6613 , n6612 );
and ( n6614 , n39 , n5429 );
or ( n6615 , n3819 , n90 );
nand ( n6616 , n6615 , n5822 );
and ( n6617 , n3609 , n6616 );
nor ( n6618 , n6614 , n6617 );
or ( n6619 , n2731 , n6613 , n5814 , n6618 );
nand ( n6620 , n6601 , n6605 , n6611 , n6619 );
nor ( n6621 , n6598 , n6600 , n6620 );
nand ( n6622 , n6589 , n6590 , n6621 );
or ( n6623 , n6491 , n6622 );
nand ( n6624 , n6623 , n4 );
nor ( n6625 , n3749 , n2636 );
nand ( n6626 , n6625 , n5823 , n3516 , n6440 );
not ( n6627 , n5831 );
nor ( n6628 , n6627 , n6441 );
nand ( n6629 , n3516 , n4166 , n40 , n6628 );
nor ( n6630 , n1 , n38 );
not ( n6631 , n6630 );
nand ( n6632 , n5 , n3516 );
nor ( n6633 , n6631 , n6344 , n6610 , n6632 );
nand ( n6634 , n6633 , n2298 , n3569 );
not ( n6635 , n4193 );
or ( n6636 , n4046 , n5852 );
and ( n6637 , n4102 , n5839 );
not ( n6638 , n17 );
and ( n6639 , n3836 , n6473 , n5827 );
and ( n6640 , n6476 , n4014 );
nor ( n6641 , n6639 , n6640 );
or ( n6642 , n6638 , n6641 );
and ( n6643 , n3836 , n3882 , n5827 );
and ( n6644 , n6482 , n4014 );
nor ( n6645 , n6643 , n6644 );
nand ( n6646 , n6642 , n6645 );
nor ( n6647 , n6637 , n6646 );
nand ( n6648 , n6636 , n6647 );
nand ( n6649 , n6635 , n4166 , n2508 , n6648 );
and ( n6650 , n6626 , n6629 , n6634 , n6649 );
nor ( n6651 , n3749 , n6464 );
and ( n6652 , n6651 , n3898 , n6440 );
not ( n6653 , n3516 );
nor ( n6654 , n4167 , n6441 );
and ( n6655 , n6339 , n6653 , n6654 );
nor ( n6656 , n6652 , n6655 );
and ( n6657 , n3281 , n4429 );
and ( n6658 , n2679 , n6365 );
nor ( n6659 , n6657 , n6658 );
not ( n6660 , n6659 );
not ( n6661 , n3276 );
not ( n6662 , n5663 );
or ( n6663 , n6661 , n6662 );
and ( n6664 , n6287 , n6358 );
not ( n6665 , n6412 );
and ( n6666 , n2467 , n3275 );
nor ( n6667 , n6666 , n6366 );
nor ( n6668 , n6664 , n6665 , n6667 );
nand ( n6669 , n6663 , n6668 );
not ( n6670 , n3265 );
not ( n6671 , n6339 );
or ( n6672 , n6670 , n6671 );
not ( n6673 , n93 );
and ( n6674 , n14 , n6673 );
not ( n6675 , n6674 );
nor ( n6676 , n841 , n6675 );
not ( n6677 , n16 );
nor ( n6678 , n19 , n2244 );
nand ( n6679 , n6677 , n6678 );
nor ( n6680 , n20 , n6679 );
or ( n6681 , n6676 , n6680 );
nand ( n6682 , n6681 , n5715 );
nand ( n6683 , n6672 , n6682 );
nor ( n6684 , n6660 , n6400 , n6669 , n6683 );
and ( n6685 , n453 , n5714 );
and ( n6686 , n5533 , n908 , n3430 );
not ( n6687 , n2493 );
and ( n6688 , n6687 , n4670 );
nor ( n6689 , n6686 , n6688 );
nand ( n6690 , n2475 , n4937 );
not ( n6691 , n3417 );
nand ( n6692 , n6691 , n4816 );
nand ( n6693 , n6689 , n6690 , n6692 );
nor ( n6694 , n6685 , n6693 );
not ( n6695 , n20 );
and ( n6696 , n6695 , n2538 , n5729 );
nor ( n6697 , n2462 , n4892 );
nor ( n6698 , n6696 , n6697 );
and ( n6699 , n6684 , n6694 , n6698 , n6422 );
not ( n6700 , n6367 );
nand ( n6701 , n2544 , n4326 );
nand ( n6702 , n6700 , n6380 , n6390 , n6701 );
or ( n6703 , n2431 , n4397 );
nand ( n6704 , n6703 , n6370 );
nor ( n6705 , n6702 , n6359 , n6704 );
and ( n6706 , n2451 , n4480 );
not ( n6707 , n2436 );
nor ( n6708 , n2501 , n4749 );
not ( n6709 , n6708 );
or ( n6710 , n6707 , n6709 );
nand ( n6711 , n4990 , n2398 , n6426 );
nand ( n6712 , n6710 , n6711 );
nor ( n6713 , n6706 , n6405 , n6712 );
and ( n6714 , n3150 , n4587 );
nor ( n6715 , n4876 , n628 , n2498 );
nor ( n6716 , n6714 , n6715 );
nand ( n6717 , n6699 , n6705 , n6713 , n6716 );
nand ( n6718 , n6355 , n2517 , n2508 , n6717 );
nand ( n6719 , n2303 , n5851 );
not ( n6720 , n6719 );
and ( n6721 , n2615 , n6720 );
not ( n6722 , n23 );
not ( n6723 , n2879 );
or ( n6724 , n6722 , n6723 , n1316 );
nor ( n6725 , n14 , n19 );
nand ( n6726 , n16 , n6725 );
or ( n6727 , n6726 , n5104 );
nand ( n6728 , n6724 , n6727 );
or ( n6729 , n1995 , n6719 );
not ( n6730 , n1407 );
not ( n6731 , n5104 );
and ( n6732 , n6730 , n6731 );
or ( n6733 , n2303 , n14 , n1929 );
or ( n6734 , n2537 , n1929 );
nand ( n6735 , n6733 , n6734 );
nor ( n6736 , n6732 , n6735 );
nand ( n6737 , n6729 , n6736 );
nor ( n6738 , n6721 , n6728 , n6737 );
or ( n6739 , n3471 , n6738 );
not ( n6740 , n18 );
not ( n6741 , n6740 );
not ( n6742 , n2868 );
not ( n6743 , n6742 );
and ( n6744 , n6741 , n6743 );
not ( n6745 , n20 );
nor ( n6746 , n6745 , n1893 );
nor ( n6747 , n6744 , n6746 );
or ( n6748 , n6747 , n6719 );
nand ( n6749 , n6739 , n6748 );
not ( n6750 , n6749 );
and ( n6751 , n5280 , n2838 , n2863 );
nor ( n6752 , n5244 , n2766 , n2843 );
nor ( n6753 , n6751 , n6752 );
and ( n6754 , n2800 , n4750 );
or ( n6755 , n2791 , n4397 );
nand ( n6756 , n2802 , n4480 );
nand ( n6757 , n6755 , n6756 );
nor ( n6758 , n6754 , n6757 );
not ( n6759 , n6758 );
and ( n6760 , n1406 , n6759 );
nor ( n6761 , n19 , n3471 );
nand ( n6762 , n16 , n6761 );
nor ( n6763 , n2766 , n6762 );
and ( n6764 , n6763 , n4670 );
nor ( n6765 , n6760 , n6764 );
or ( n6766 , n2488 , n5275 );
nand ( n6767 , n6766 , n6383 );
and ( n6768 , n18 , n6767 );
not ( n6769 , n2800 );
not ( n6770 , n5282 );
or ( n6771 , n6769 , n6770 );
and ( n6772 , n5167 , n2538 , n5292 );
nor ( n6773 , n6772 , n6381 );
nand ( n6774 , n6771 , n6773 );
and ( n6775 , n1582 , n6774 );
nor ( n6776 , n6768 , n6775 );
not ( n6777 , n23 );
not ( n6778 , n2781 );
or ( n6779 , n6777 , n20 , n6778 );
nand ( n6780 , n6779 , n2971 );
and ( n6781 , n6780 , n18 , n5270 );
not ( n6782 , n2879 );
nor ( n6783 , n6782 , n1316 , n5248 , n308 );
nor ( n6784 , n6781 , n6783 );
and ( n6785 , n6753 , n6765 , n6776 , n6784 );
or ( n6786 , n6006 , n2791 , n4417 );
or ( n6787 , n5284 , n2450 , n5286 );
nand ( n6788 , n6786 , n6787 );
and ( n6789 , n309 , n6788 );
or ( n6790 , n2228 , n6719 );
not ( n6791 , n14 );
not ( n6792 , n2744 );
not ( n6793 , n1891 );
not ( n6794 , n6793 );
or ( n6795 , n6792 , n6794 );
nand ( n6796 , n6795 , n23 );
or ( n6797 , n6791 , n6796 );
nand ( n6798 , n6790 , n6797 );
and ( n6799 , n2066 , n6798 );
not ( n6800 , n18 );
or ( n6801 , n6800 , n6738 );
nand ( n6802 , n16 , n1554 , n6798 );
nand ( n6803 , n6801 , n6802 );
nor ( n6804 , n6789 , n6799 , n6803 );
not ( n6805 , n1891 );
nor ( n6806 , n6805 , n912 );
or ( n6807 , n2543 , n6806 );
nand ( n6808 , n6807 , n23 );
not ( n6809 , n18 );
or ( n6810 , n5035 , n2488 );
nand ( n6811 , n6810 , n6701 );
nand ( n6812 , n6809 , n6811 );
not ( n6813 , n18 );
not ( n6814 , n4585 );
or ( n6815 , n6814 , n2745 );
or ( n6816 , n14 , n6796 );
nand ( n6817 , n6815 , n6816 );
and ( n6818 , n454 , n6817 );
and ( n6819 , n2538 , n4427 );
and ( n6820 , n2802 , n5663 );
nor ( n6821 , n6819 , n6820 );
nor ( n6822 , n20 , n6821 );
nor ( n6823 , n6818 , n6822 );
not ( n6824 , n20 );
and ( n6825 , n6824 , n6737 );
and ( n6826 , n6742 , n6286 , n455 );
nor ( n6827 , n6826 , n6719 );
nor ( n6828 , n6825 , n6827 );
and ( n6829 , n4940 , n6780 );
not ( n6830 , n20 );
or ( n6831 , n2789 , n4815 );
and ( n6832 , n23 , n2879 , n96 );
not ( n6833 , n3298 );
nand ( n6834 , n16 , n6833 );
not ( n6835 , n6834 );
and ( n6836 , n6835 , n5149 );
nor ( n6837 , n6832 , n6836 );
nand ( n6838 , n6831 , n6837 );
and ( n6839 , n6830 , n6838 );
nor ( n6840 , n6829 , n6839 );
nand ( n6841 , n6823 , n6828 , n6840 );
nand ( n6842 , n6813 , n6841 );
and ( n6843 , n6808 , n6812 , n6842 );
nand ( n6844 , n6750 , n6785 , n6804 , n6843 );
nand ( n6845 , n6355 , n1971 , n2508 , n6844 );
and ( n6846 , n6650 , n6656 , n6718 , n6845 );
not ( n6847 , n6628 );
nor ( n6848 , n6847 , n6632 );
and ( n6849 , n6848 , n3569 , n445 );
nand ( n6850 , n4166 , n2507 , n38 , n3531 );
not ( n6851 , n6654 );
and ( n6852 , n6850 , n6851 );
nor ( n6853 , n6852 , n6442 );
nor ( n6854 , n6849 , n6853 );
not ( n6855 , n2507 );
nor ( n6856 , n6338 , n4082 , n6855 );
nor ( n6857 , n3516 , n3749 );
and ( n6858 , n6856 , n6857 , n3531 );
not ( n6859 , n6857 );
nand ( n6860 , n2507 , n4013 );
nor ( n6861 , n6859 , n6344 , n6464 , n6860 );
nor ( n6862 , n6858 , n6861 );
and ( n6863 , n6846 , n6854 , n6862 );
not ( n6864 , n3371 );
and ( n6865 , n6757 , n1406 , n6864 );
and ( n6866 , n16 , n5410 );
or ( n6867 , n5868 , n42 );
or ( n6868 , n2303 , n5409 );
nand ( n6869 , n6867 , n6868 );
nand ( n6870 , n3331 , n6869 );
not ( n6871 , n6870 );
nor ( n6872 , n6866 , n6871 );
not ( n6873 , n2438 );
nor ( n6874 , n6872 , n6873 , n2182 );
nor ( n6875 , n6865 , n6874 );
not ( n6876 , n6875 );
not ( n6877 , n5533 );
nand ( n6878 , n908 , n2183 );
or ( n6879 , n6877 , n2498 , n6878 );
and ( n6880 , n3352 , n6869 );
not ( n6881 , n16 );
and ( n6882 , n6881 , n5410 );
nor ( n6883 , n6880 , n6882 );
or ( n6884 , n6878 , n6883 );
nand ( n6885 , n6879 , n6884 );
and ( n6886 , n435 , n6869 );
and ( n6887 , n2332 , n5410 );
nor ( n6888 , n6886 , n6887 );
or ( n6889 , n6888 , n3471 , n3371 );
not ( n6890 , n4671 );
nand ( n6891 , n6890 , n1314 , n3428 );
nand ( n6892 , n6889 , n6891 );
or ( n6893 , n3371 , n1415 , n6870 );
not ( n6894 , n5410 );
not ( n6895 , n1921 );
or ( n6896 , n6894 , n6895 , n3371 );
nand ( n6897 , n6893 , n6896 );
nor ( n6898 , n6876 , n6885 , n6892 , n6897 );
and ( n6899 , n782 , n6869 );
nand ( n6900 , n3345 , n5410 );
nand ( n6901 , n6900 , n6701 );
nor ( n6902 , n6899 , n6901 );
not ( n6903 , n2192 );
not ( n6904 , n6883 );
and ( n6905 , n6903 , n6904 );
nor ( n6906 , n6905 , n6697 , n6822 );
and ( n6907 , n3413 , n5653 );
or ( n6908 , n841 , n6872 );
nand ( n6909 , n6908 , n6692 );
nor ( n6910 , n6907 , n6909 );
not ( n6911 , n20 );
not ( n6912 , n6888 );
and ( n6913 , n6911 , n6912 );
not ( n6914 , n3025 );
nor ( n6915 , n6914 , n4586 );
nor ( n6916 , n6913 , n6915 , n6715 );
nand ( n6917 , n6902 , n6906 , n6910 , n6916 );
and ( n6918 , n2183 , n6917 );
nand ( n6919 , n1730 , n5798 , n2736 , n4990 );
nand ( n6920 , n6708 , n1314 , n5798 );
nand ( n6921 , n6919 , n6920 );
and ( n6922 , n570 , n6869 );
and ( n6923 , n1919 , n5410 );
not ( n6924 , n19 );
or ( n6925 , n6924 , n6883 );
nand ( n6926 , n6925 , n6900 );
nor ( n6927 , n6922 , n6923 , n6926 );
and ( n6928 , n2559 , n5280 );
and ( n6929 , n942 , n6869 );
nor ( n6930 , n6928 , n6929 );
nand ( n6931 , n2544 , n4319 );
nand ( n6932 , n6927 , n6930 , n6931 , n6378 );
not ( n6933 , n6932 );
and ( n6934 , n3413 , n5262 );
not ( n6935 , n6376 );
and ( n6936 , n2489 , n5482 );
nor ( n6937 , n3417 , n5244 );
nor ( n6938 , n6936 , n6937 );
not ( n6939 , n20 );
nand ( n6940 , n6939 , n6788 );
nand ( n6941 , n6935 , n6938 , n6940 );
not ( n6942 , n6428 );
nand ( n6943 , n6395 , n6942 );
nor ( n6944 , n6934 , n6941 , n6943 );
not ( n6945 , n19 );
not ( n6946 , n6872 );
and ( n6947 , n6945 , n6946 );
not ( n6948 , n20 );
nor ( n6949 , n6948 , n6773 );
nor ( n6950 , n6947 , n6949 );
nand ( n6951 , n6944 , n6950 , n6888 , n6421 );
not ( n6952 , n6951 );
and ( n6953 , n6933 , n6952 );
nor ( n6954 , n6953 , n3440 );
nor ( n6955 , n6918 , n6921 , n6954 );
not ( n6956 , n3228 );
not ( n6957 , n6701 );
and ( n6958 , n6956 , n6957 );
not ( n6959 , n13 );
nand ( n6960 , n6959 , n1406 );
not ( n6961 , n6960 );
or ( n6962 , n2306 , n6244 );
nor ( n6963 , n5575 , n5572 );
or ( n6964 , n1407 , n6963 );
nand ( n6965 , n42 , n5429 );
or ( n6966 , n795 , n6965 );
nand ( n6967 , n6962 , n6964 , n6966 );
and ( n6968 , n6961 , n6967 );
nor ( n6969 , n6958 , n6968 );
not ( n6970 , n6969 );
not ( n6971 , n19 );
nor ( n6972 , n6971 , n6960 );
not ( n6973 , n6972 );
or ( n6974 , n6244 , n42 );
nand ( n6975 , n6974 , n6965 );
not ( n6976 , n6975 );
or ( n6977 , n6976 , n521 );
or ( n6978 , n16 , n6963 );
nand ( n6979 , n6977 , n6978 );
not ( n6980 , n6979 );
or ( n6981 , n6973 , n6980 );
not ( n6982 , n13 );
not ( n6983 , n19 );
nor ( n6984 , n2234 , n3471 );
or ( n6985 , n2396 , n6244 );
and ( n6986 , n2398 , n5429 );
and ( n6987 , n17 , n5873 );
nor ( n6988 , n6986 , n6987 );
nand ( n6989 , n6985 , n6988 );
nand ( n6990 , n6982 , n6983 , n6984 , n6989 );
nand ( n6991 , n6981 , n6990 );
or ( n6992 , n4397 , n6960 , n3309 );
and ( n6993 , n6961 , n3299 );
nor ( n6994 , n1415 , n3247 );
nor ( n6995 , n6993 , n6994 );
not ( n6996 , n6989 );
or ( n6997 , n6995 , n6996 );
nand ( n6998 , n6992 , n6997 );
nand ( n6999 , n1924 , n6975 );
or ( n7000 , n13 , n6999 );
not ( n7001 , n13 );
nand ( n7002 , n5103 , n1921 , n7001 , n5429 );
nand ( n7003 , n7000 , n7002 );
nor ( n7004 , n6970 , n6991 , n6998 , n7003 );
nor ( n7005 , n2437 , n3228 );
and ( n7006 , n7005 , n6708 );
and ( n7007 , n724 , n6975 );
not ( n7008 , n6963 );
and ( n7009 , n16 , n7008 );
nor ( n7010 , n7007 , n7009 );
or ( n7011 , n7010 , n2437 , n3228 );
or ( n7012 , n6960 , n6756 );
nand ( n7013 , n7011 , n7012 );
and ( n7014 , n942 , n6975 );
or ( n7015 , n2433 , n7010 );
and ( n7016 , n20 , n6967 );
and ( n7017 , n908 , n6979 );
nor ( n7018 , n7016 , n7017 );
nand ( n7019 , n7015 , n7018 );
nand ( n7020 , n6382 , n6395 );
nor ( n7021 , n7014 , n7019 , n7020 );
and ( n7022 , n6369 , n6989 );
nor ( n7023 , n5430 , n5405 , n1920 );
nor ( n7024 , n7022 , n7023 , n6372 );
and ( n7025 , n2389 , n6989 );
nor ( n7026 , n7025 , n6392 );
and ( n7027 , n7026 , n6931 , n6429 );
and ( n7028 , n7021 , n7024 , n7027 );
nor ( n7029 , n7028 , n3236 );
nor ( n7030 , n7006 , n7013 , n7029 );
not ( n7031 , n19 );
and ( n7032 , n7031 , n2398 , n6984 );
not ( n7033 , n13 );
and ( n7034 , n7032 , n7033 , n6890 );
and ( n7035 , n5533 , n6972 , n3430 );
nor ( n7036 , n7034 , n7035 );
and ( n7037 , n766 , n6975 );
nand ( n7038 , n17 , n3246 );
not ( n7039 , n7038 );
and ( n7040 , n5873 , n624 , n7039 );
not ( n7041 , n20 );
not ( n7042 , n16 );
and ( n7043 , n7041 , n7042 , n5575 );
nor ( n7044 , n7040 , n7043 );
not ( n7045 , n7044 );
nor ( n7046 , n20 , n2791 , n5430 );
nor ( n7047 , n7037 , n7045 , n7046 );
and ( n7048 , n3278 , n6989 );
and ( n7049 , n6680 , n5873 );
nor ( n7050 , n7048 , n7049 );
or ( n7051 , n2243 , n2515 );
nand ( n7052 , n7051 , n6989 );
and ( n7053 , n7047 , n7050 , n6378 , n7052 );
and ( n7054 , n3265 , n6245 );
or ( n7055 , n2443 , n3128 , n6419 );
nand ( n7056 , n5285 , n3276 , n5289 );
nand ( n7057 , n7055 , n7056 );
nor ( n7058 , n841 , n7010 );
nor ( n7059 , n7054 , n7057 , n7058 );
and ( n7060 , n570 , n6975 );
nor ( n7061 , n6006 , n3270 , n5258 );
nor ( n7062 , n5430 , n5405 , n3346 );
nor ( n7063 , n7060 , n7061 , n7062 );
nor ( n7064 , n3407 , n632 );
and ( n7065 , n7064 , n5262 );
nor ( n7066 , n7065 , n6415 , n6376 );
nand ( n7067 , n7053 , n7059 , n7063 , n7066 );
and ( n7068 , n3250 , n7067 );
and ( n7069 , n782 , n6975 );
or ( n7070 , n2242 , n6996 );
or ( n7071 , n3408 , n4892 );
nand ( n7072 , n7070 , n7071 );
nor ( n7073 , n7069 , n7072 , n7062 );
and ( n7074 , n2468 , n6989 );
and ( n7075 , n2447 , n4429 );
and ( n7076 , n2418 , n5663 );
nor ( n7077 , n7074 , n7075 , n7076 );
not ( n7078 , n20 );
and ( n7079 , n7078 , n6967 );
nor ( n7080 , n7079 , n6915 , n6715 );
and ( n7081 , n2478 , n4816 );
and ( n7082 , n629 , n6979 );
nor ( n7083 , n7081 , n7082 );
not ( n7084 , n7058 );
and ( n7085 , n7083 , n7084 , n6690 );
nand ( n7086 , n7073 , n7077 , n7080 , n7085 );
and ( n7087 , n3121 , n7086 );
not ( n7088 , n6994 );
nor ( n7089 , n2443 , n7088 );
and ( n7090 , n7089 , n4990 );
nor ( n7091 , n7068 , n7087 , n7090 );
nand ( n7092 , n7004 , n7030 , n7036 , n7091 );
and ( n7093 , n3119 , n7092 );
and ( n7094 , n994 , n6844 );
nor ( n7095 , n7093 , n7094 );
not ( n7096 , n2 );
nand ( n7097 , n1849 , n6844 );
not ( n7098 , n6137 );
nand ( n7099 , n7098 , n2998 , n2517 );
and ( n7100 , n454 , n2938 );
and ( n7101 , n7100 , n5984 );
or ( n7102 , n5248 , n2186 , n2745 );
nand ( n7103 , n7102 , n6940 );
nor ( n7104 , n7101 , n7103 , n6937 );
not ( n7105 , n2678 );
not ( n7106 , n6796 );
and ( n7107 , n7105 , n7106 );
and ( n7108 , n6837 , n6736 );
nor ( n7109 , n7108 , n20 );
nor ( n7110 , n7107 , n7109 );
nand ( n7111 , n2461 , n5270 );
or ( n7112 , n6014 , n6275 );
nand ( n7113 , n7112 , n2998 );
nand ( n7114 , n7104 , n7110 , n7111 , n7113 );
and ( n7115 , n1982 , n7114 );
and ( n7116 , n3069 , n6774 );
nor ( n7117 , n7115 , n7116 );
nand ( n7118 , n7099 , n7117 );
or ( n7119 , n3549 , n6821 );
not ( n7120 , n3035 );
and ( n7121 , n6064 , n2066 , n7120 );
and ( n7122 , n3070 , n3549 );
nor ( n7123 , n7122 , n6736 );
nor ( n7124 , n7121 , n7123 );
nand ( n7125 , n7119 , n7124 );
and ( n7126 , n3069 , n6728 );
or ( n7127 , n6797 , n3079 );
or ( n7128 , n2579 , n6808 );
nand ( n7129 , n7127 , n7128 );
and ( n7130 , n3435 , n3074 , n2303 , n5959 );
nor ( n7131 , n7126 , n7129 , n7130 );
and ( n7132 , n5280 , n2838 , n3080 );
and ( n7133 , n3056 , n5943 );
nor ( n7134 , n7132 , n7133 );
not ( n7135 , n3549 );
nand ( n7136 , n6817 , n2816 , n7135 );
nand ( n7137 , n454 , n2517 , n2938 , n6096 );
nand ( n7138 , n7131 , n7134 , n7136 , n7137 );
nor ( n7139 , n7118 , n7125 , n7138 );
and ( n7140 , n2954 , n6198 );
not ( n7141 , n20 );
or ( n7142 , n7141 , n6758 );
or ( n7143 , n2067 , n6797 );
nand ( n7144 , n7142 , n7143 , n6808 );
nor ( n7145 , n7140 , n7144 , n6811 );
not ( n7146 , n6736 );
or ( n7147 , n6728 , n7146 );
nand ( n7148 , n7147 , n20 );
nand ( n7149 , n6890 , n2066 , n2838 );
not ( n7150 , n6311 );
and ( n7151 , n7150 , n2066 , n2977 );
and ( n7152 , n2303 , n6260 );
nor ( n7153 , n7151 , n7152 );
nand ( n7154 , n7145 , n7148 , n7149 , n7153 );
nand ( n7155 , n2517 , n7154 );
and ( n7156 , n6294 , n2998 , n2517 );
not ( n7157 , n6838 );
or ( n7158 , n3549 , n7157 );
and ( n7159 , n6266 , n2920 , n1982 );
and ( n7160 , n1982 , n6767 );
nor ( n7161 , n7159 , n7160 );
nand ( n7162 , n4940 , n2461 , n2517 );
nand ( n7163 , n7158 , n7161 , n7162 );
nor ( n7164 , n7156 , n7163 );
nand ( n7165 , n7097 , n7139 , n7155 , n7164 );
nand ( n7166 , n7096 , n7165 );
nand ( n7167 , n6898 , n6955 , n7095 , n7166 );
nand ( n7168 , n7167 , n2506 , n4254 );
not ( n7169 , n4151 );
or ( n7170 , n6618 , n5814 , n6445 );
nand ( n7171 , n3516 , n4081 );
not ( n7172 , n3372 );
or ( n7173 , n7171 , n7172 , n5809 );
nand ( n7174 , n7170 , n7173 );
not ( n7175 , n5800 );
or ( n7176 , n3373 , n4082 , n7175 );
and ( n7177 , n994 , n6648 );
and ( n7178 , n38 , n5869 );
nor ( n7179 , n7177 , n7178 );
nand ( n7180 , n7176 , n7179 );
nor ( n7181 , n7174 , n7180 );
and ( n7182 , n3836 , n5862 , n6454 );
and ( n7183 , n5844 , n4082 , n3119 );
nor ( n7184 , n7182 , n7183 );
not ( n7185 , n5874 );
not ( n7186 , n13 );
nand ( n7187 , n7185 , n7186 , n6612 );
not ( n7188 , n2 );
not ( n7189 , n6041 );
nand ( n7190 , n7189 , n6061 );
nand ( n7191 , n7190 , n4051 , n1982 );
and ( n7192 , n4056 , n6158 );
and ( n7193 , n2649 , n6646 );
not ( n7194 , n6641 );
and ( n7195 , n2245 , n7194 );
not ( n7196 , n6645 );
and ( n7197 , n14 , n7196 );
nor ( n7198 , n7195 , n7197 );
or ( n7199 , n2067 , n7198 );
not ( n7200 , n6646 );
or ( n7201 , n912 , n7200 );
nand ( n7202 , n7199 , n7201 );
nor ( n7203 , n7192 , n7193 , n7202 );
not ( n7204 , n4054 );
not ( n7205 , n7204 );
not ( n7206 , n6162 );
and ( n7207 , n7205 , n7206 );
and ( n7208 , n4048 , n6226 );
nor ( n7209 , n7207 , n7208 );
not ( n7210 , n4047 );
not ( n7211 , n6555 );
or ( n7212 , n7210 , n7211 );
not ( n7213 , n4059 );
nand ( n7214 , n7213 , n6191 );
nand ( n7215 , n7212 , n7214 );
not ( n7216 , n7215 );
nand ( n7217 , n7203 , n7209 , n7216 );
nand ( n7218 , n7217 , n2517 );
not ( n7219 , n4048 );
not ( n7220 , n6152 );
or ( n7221 , n7219 , n7220 );
not ( n7222 , n4091 );
and ( n7223 , n7222 , n6126 );
not ( n7224 , n4047 );
not ( n7225 , n6144 );
or ( n7226 , n7224 , n7225 );
nand ( n7227 , n4020 , n6122 );
nand ( n7228 , n7226 , n7227 );
nor ( n7229 , n7223 , n7228 );
nand ( n7230 , n4093 , n6133 );
nand ( n7231 , n7221 , n7229 , n7230 );
or ( n7232 , n2186 , n7198 );
and ( n7233 , n6096 , n4020 , n2615 );
and ( n7234 , n4085 , n6129 );
nor ( n7235 , n7233 , n7234 );
or ( n7236 , n2189 , n4134 );
nand ( n7237 , n7236 , n6646 );
nand ( n7238 , n7232 , n7235 , n7237 );
or ( n7239 , n7231 , n7238 );
nand ( n7240 , n7239 , n2517 );
and ( n7241 , n7191 , n7218 , n7240 );
or ( n7242 , n2579 , n4048 , n5976 );
and ( n7243 , n5940 , n4060 , n1982 );
and ( n7244 , n5943 , n4047 , n3069 );
nor ( n7245 , n7243 , n7244 );
nand ( n7246 , n7242 , n7245 );
nand ( n7247 , n4048 , n3080 );
or ( n7248 , n7247 , n2228 , n6074 );
or ( n7249 , n6068 , n4048 , n2602 );
nand ( n7250 , n7248 , n7249 );
nand ( n7251 , n450 , n2816 , n1982 );
or ( n7252 , n5989 , n4091 , n7251 );
nand ( n7253 , n6518 , n6018 );
or ( n7254 , n7253 , n38 );
nand ( n7255 , n7252 , n7254 );
nor ( n7256 , n7246 , n7250 , n7255 );
not ( n7257 , n4081 );
nand ( n7258 , n7257 , n3080 , n2229 , n6064 );
and ( n7259 , n1849 , n6648 );
and ( n7260 , n3074 , n6646 );
nor ( n7261 , n7259 , n7260 );
and ( n7262 , n6646 , n4074 , n3069 );
not ( n7263 , n4020 );
nor ( n7264 , n6043 , n7263 , n7251 );
nor ( n7265 , n7262 , n7264 );
nand ( n7266 , n7261 , n7265 );
or ( n7267 , n6641 , n3789 , n6493 );
or ( n7268 , n6645 , n2579 , n2678 );
nand ( n7269 , n7267 , n7268 );
or ( n7270 , n3079 , n7198 );
or ( n7271 , n6529 , n6509 );
nand ( n7272 , n7271 , n6646 );
nand ( n7273 , n7270 , n7272 );
nor ( n7274 , n7266 , n7269 , n7273 );
nand ( n7275 , n7241 , n7256 , n7258 , n7274 );
and ( n7276 , n7188 , n7275 );
not ( n7277 , n3119 );
nor ( n7278 , n7277 , n4081 , n5836 , n6246 );
nor ( n7279 , n7276 , n7278 );
nand ( n7280 , n7181 , n7184 , n7187 , n7279 );
nand ( n7281 , n7169 , n7280 );
and ( n7282 , n6863 , n7168 , n7281 );
nand ( n7283 , n6436 , n6624 , n7282 );
and ( n7284 , n4238 , n7283 );
nor ( n7285 , n5310 , n7284 );
not ( n7286 , n4267 );
nand ( n7287 , n7286 , n6844 );
and ( n7288 , n4244 , n6330 );
and ( n7289 , n23 , n4263 );
nor ( n7290 , n7288 , n7289 );
and ( n7291 , n4277 , n7165 );
and ( n7292 , n4271 , n5239 );
and ( n7293 , n4259 , n6315 );
nor ( n7294 , n7291 , n7292 , n7293 );
nand ( n7295 , n7285 , n7287 , n7290 , n7294 );
nor ( n7296 , n4261 , n4240 );
not ( n7297 , n24 );
not ( n7298 , n34 );
not ( n7299 , n7298 );
not ( n7300 , n190 );
nor ( n7301 , n7300 , n30 );
not ( n7302 , n7301 );
not ( n7303 , n7302 );
not ( n7304 , n45 );
not ( n7305 , n133 );
or ( n7306 , n7304 , n7305 );
nand ( n7307 , n28 , n44 );
nand ( n7308 , n7306 , n7307 );
buf ( n7309 , n7308 );
nand ( n7310 , n7303 , n7309 );
nand ( n7311 , n166 , n30 );
not ( n7312 , n7311 );
not ( n7313 , n171 );
not ( n7314 , n45 );
nand ( n7315 , n27 , n7314 );
not ( n7316 , n7315 );
or ( n7317 , n7313 , n7316 );
nand ( n7318 , n7317 , n7307 );
nand ( n7319 , n7312 , n7318 );
not ( n7320 , n191 );
not ( n7321 , n189 );
or ( n7322 , n7320 , n7321 );
nand ( n7323 , n191 , n36 );
nand ( n7324 , n7322 , n7323 );
and ( n7325 , n7308 , n7324 );
nor ( n7326 , n7323 , n4353 );
nor ( n7327 , n7325 , n7326 );
buf ( n7328 , n7327 );
nand ( n7329 , n7310 , n7319 , n7328 );
not ( n7330 , n7329 );
or ( n7331 , n7299 , n7330 );
not ( n7332 , n4404 );
buf ( n7333 , n7332 );
not ( n7334 , n7333 );
not ( n7335 , n7312 );
and ( n7336 , n7334 , n7335 );
buf ( n7337 , n7318 );
not ( n7338 , n7337 );
nor ( n7339 , n7336 , n7338 );
not ( n7340 , n7328 );
or ( n7341 , n7339 , n7340 );
or ( n7342 , n30 , n34 );
nand ( n7343 , n7341 , n7342 );
nand ( n7344 , n7331 , n7343 );
not ( n7345 , n7344 );
not ( n7346 , n7345 );
and ( n7347 , n25 , n7346 );
nand ( n7348 , n221 , n4306 );
not ( n7349 , n7309 );
and ( n7350 , n7348 , n7349 );
nor ( n7351 , n7350 , n2317 );
not ( n7352 , n7351 );
not ( n7353 , n350 );
nand ( n7354 , n7333 , n7309 );
not ( n7355 , n7309 );
nor ( n7356 , n7335 , n7355 );
and ( n7357 , n7319 , n7327 );
nor ( n7358 , n7357 , n30 );
nor ( n7359 , n7356 , n7358 );
and ( n7360 , n7354 , n7359 );
not ( n7361 , n7360 );
nand ( n7362 , n7353 , n7361 );
nand ( n7363 , n7352 , n7362 );
nor ( n7364 , n7347 , n7363 );
or ( n7365 , n7297 , n7364 );
not ( n7366 , n24 );
nor ( n7367 , n7366 , n4315 );
not ( n7368 , n7367 );
not ( n7369 , n2317 );
not ( n7370 , n7369 );
not ( n7371 , n7370 );
or ( n7372 , n7371 , n7360 );
nand ( n7373 , n7372 , n7352 );
not ( n7374 , n4311 );
nand ( n7375 , n7373 , n7374 , n3604 );
nand ( n7376 , n7368 , n7375 );
not ( n7377 , n7376 );
nand ( n7378 , n7365 , n7377 );
nand ( n7379 , n3800 , n18 , n3521 );
not ( n7380 , n7379 );
and ( n7381 , n7378 , n7380 , n2463 );
and ( n7382 , n998 , n7374 );
buf ( n7383 , n2317 );
not ( n7384 , n7383 );
nand ( n7385 , n7333 , n7337 );
nand ( n7386 , n7385 , n7319 , n7328 );
not ( n7387 , n7386 );
or ( n7388 , n7384 , n7387 );
nand ( n7389 , n7388 , n7352 );
nand ( n7390 , n24 , n7382 , n7389 );
not ( n7391 , n24 );
and ( n7392 , n7391 , n7382 , n7373 );
nand ( n7393 , n24 , n111 );
not ( n7394 , n7393 );
nor ( n7395 , n7392 , n7394 );
nand ( n7396 , n7390 , n7395 );
and ( n7397 , n2303 , n450 , n7396 );
not ( n7398 , n14 );
not ( n7399 , n17 );
not ( n7400 , n7349 );
nand ( n7401 , n7382 , n7400 );
and ( n7402 , n7393 , n7401 );
nor ( n7403 , n7402 , n15 );
not ( n7404 , n7403 );
or ( n7405 , n7399 , n7404 );
not ( n7406 , n7393 );
not ( n7407 , n7307 );
nand ( n7408 , n7407 , n7382 );
not ( n7409 , n7408 );
or ( n7410 , n7406 , n7409 );
not ( n7411 , n17 );
nand ( n7412 , n7410 , n7411 );
nand ( n7413 , n7405 , n7412 );
nand ( n7414 , n7398 , n7413 );
not ( n7415 , n7414 );
nor ( n7416 , n7397 , n7415 );
nor ( n7417 , n3089 , n7416 );
and ( n7418 , n7380 , n7417 );
nor ( n7419 , n7381 , n7418 );
not ( n7420 , n24 );
not ( n7421 , n25 );
not ( n7422 , n7337 );
and ( n7423 , n7422 , n7328 );
nor ( n7424 , n7423 , n391 );
nor ( n7425 , n7424 , n7329 );
not ( n7426 , n7425 );
not ( n7427 , n7426 );
not ( n7428 , n7427 );
not ( n7429 , n7428 );
not ( n7430 , n7429 );
not ( n7431 , n7430 );
or ( n7432 , n7421 , n7431 );
not ( n7433 , n7363 );
nand ( n7434 , n7432 , n7433 );
not ( n7435 , n7434 );
or ( n7436 , n7420 , n7435 );
nand ( n7437 , n7436 , n7377 );
and ( n7438 , n7437 , n7380 , n2544 );
not ( n7439 , n554 );
not ( n7440 , n7439 );
not ( n7441 , n7440 );
not ( n7442 , n1481 );
not ( n7443 , n7425 );
not ( n7444 , n7303 );
not ( n7445 , n7444 );
not ( n7446 , n7445 );
nand ( n7447 , n7335 , n7446 );
not ( n7448 , n4617 );
not ( n7449 , n7448 );
not ( n7450 , n7449 );
not ( n7451 , n7450 );
nand ( n7452 , n7443 , n7447 , n7451 );
nand ( n7453 , n34 , n7386 );
not ( n7454 , n7453 );
not ( n7455 , n7445 );
not ( n7456 , n7455 );
not ( n7457 , n34 );
nand ( n7458 , n7457 , n30 , n7337 );
not ( n7459 , n34 );
nand ( n7460 , n36 , n7459 , n7337 );
not ( n7461 , n7460 );
not ( n7462 , n34 );
nand ( n7463 , n7462 , n392 , n7309 );
not ( n7464 , n7463 );
or ( n7465 , n7461 , n7464 );
nand ( n7466 , n7465 , n391 );
nand ( n7467 , n7458 , n7466 );
not ( n7468 , n7467 );
or ( n7469 , n7456 , n7468 );
and ( n7470 , n391 , n7444 );
nor ( n7471 , n7470 , n385 );
nand ( n7472 , n7471 , n7386 );
nand ( n7473 , n7469 , n7472 );
nor ( n7474 , n7454 , n7473 );
nand ( n7475 , n7452 , n7474 );
not ( n7476 , n7475 );
or ( n7477 , n7442 , n7476 );
nand ( n7478 , n487 , n7344 );
nand ( n7479 , n7477 , n7478 );
or ( n7480 , n7363 , n7479 );
not ( n7481 , n7480 );
or ( n7482 , n7441 , n7481 );
not ( n7483 , n35 );
and ( n7484 , n33 , n7352 );
nand ( n7485 , n477 , n7361 );
nand ( n7486 , n7484 , n7485 );
not ( n7487 , n7486 );
not ( n7488 , n32 );
nand ( n7489 , n7488 , n7351 );
not ( n7490 , n26 );
not ( n7491 , n606 );
not ( n7492 , n7491 );
and ( n7493 , n7490 , n7492 );
nand ( n7494 , n234 , n7493 , n7361 );
nand ( n7495 , n7489 , n7494 );
not ( n7496 , n7495 );
nand ( n7497 , n382 , n7475 );
nand ( n7498 , n7496 , n7497 );
not ( n7499 , n7498 );
or ( n7500 , n7487 , n7499 );
not ( n7501 , n895 );
not ( n7502 , n7346 );
not ( n7503 , n7502 );
and ( n7504 , n7501 , n7503 );
not ( n7505 , n32 );
and ( n7506 , n7505 , n7479 );
nor ( n7507 , n7504 , n7506 );
nand ( n7508 , n7500 , n7507 );
nand ( n7509 , n7483 , n7508 );
nand ( n7510 , n7482 , n7509 );
not ( n7511 , n7510 );
not ( n7512 , n24 );
or ( n7513 , n7511 , n7512 );
nand ( n7514 , n7513 , n7377 );
not ( n7515 , n7514 );
nand ( n7516 , n2458 , n3082 );
nor ( n7517 , n7515 , n7379 , n7516 );
nor ( n7518 , n7438 , n7517 );
nor ( n7519 , n1582 , n7379 );
not ( n7520 , n24 );
not ( n7521 , n7353 );
not ( n7522 , n7521 );
not ( n7523 , n32 );
not ( n7524 , n2317 );
or ( n7525 , n7523 , n7524 );
not ( n7526 , n7525 );
not ( n7527 , n7467 );
nand ( n7528 , n7527 , n7453 );
nand ( n7529 , n7526 , n7528 );
and ( n7530 , n32 , n7351 );
not ( n7531 , n7530 );
nand ( n7532 , n236 , n7528 );
not ( n7533 , n4372 );
nor ( n7534 , n26 , n7533 );
nand ( n7535 , n234 , n7534 , n7361 );
nand ( n7536 , n7532 , n7489 , n7535 );
not ( n7537 , n7536 );
and ( n7538 , n7529 , n7531 , n7537 );
or ( n7539 , n7522 , n7538 );
nand ( n7540 , n234 , n1382 , n7361 );
and ( n7541 , n7489 , n7540 );
and ( n7542 , n7541 , n7532 );
nand ( n7543 , n7539 , n7542 , n7535 );
not ( n7544 , n7543 );
or ( n7545 , n7520 , n7544 );
nand ( n7546 , n7545 , n7377 );
and ( n7547 , n7519 , n2538 , n7546 );
nand ( n7548 , n7382 , n7337 );
and ( n7549 , n7393 , n7548 );
nor ( n7550 , n7549 , n15 );
nand ( n7551 , n17 , n7550 );
not ( n7552 , n17 );
nand ( n7553 , n7552 , n171 , n4315 );
and ( n7554 , n7553 , n7412 );
nand ( n7555 , n7551 , n7554 );
nand ( n7556 , n14 , n7555 );
nand ( n7557 , n7414 , n7556 );
not ( n7558 , n7557 );
nor ( n7559 , n19 , n7558 );
not ( n7560 , n7396 );
not ( n7561 , n17 );
nor ( n7562 , n7560 , n7561 , n19 , n2937 );
or ( n7563 , n7559 , n7562 );
and ( n7564 , n7380 , n7563 );
nor ( n7565 , n7547 , n7564 );
not ( n7566 , n24 );
not ( n7567 , n487 );
not ( n7568 , n7528 );
or ( n7569 , n7567 , n7568 );
nand ( n7570 , n534 , n7344 );
nand ( n7571 , n7569 , n7570 );
nand ( n7572 , n256 , n7571 );
nand ( n7573 , n256 , n7363 );
not ( n7574 , n33 );
and ( n7575 , n7574 , n7352 );
not ( n7576 , n222 );
not ( n7577 , n7576 );
nand ( n7578 , n7577 , n7361 );
nand ( n7579 , n7575 , n7578 );
not ( n7580 , n7579 );
not ( n7581 , n7536 );
or ( n7582 , n7580 , n7581 );
not ( n7583 , n215 );
not ( n7584 , n7345 );
and ( n7585 , n7583 , n7584 );
not ( n7586 , n32 );
and ( n7587 , n7586 , n7571 );
nor ( n7588 , n7585 , n7587 );
nand ( n7589 , n7582 , n7588 );
nand ( n7590 , n35 , n7589 );
nand ( n7591 , n7572 , n7573 , n7590 );
not ( n7592 , n7591 );
or ( n7593 , n7566 , n7592 );
nand ( n7594 , n7593 , n7377 );
nand ( n7595 , n96 , n7594 );
nand ( n7596 , n16 , n7557 );
not ( n7597 , n24 );
not ( n7598 , n1151 );
not ( n7599 , n7598 );
not ( n7600 , n7599 );
not ( n7601 , n7600 );
not ( n7602 , n7475 );
or ( n7603 , n7601 , n7602 );
nand ( n7604 , n7603 , n7570 );
or ( n7605 , n7363 , n7604 );
nand ( n7606 , n7605 , n256 );
nand ( n7607 , n7575 , n7485 );
not ( n7608 , n7607 );
not ( n7609 , n7498 );
or ( n7610 , n7608 , n7609 );
not ( n7611 , n738 );
not ( n7612 , n7502 );
and ( n7613 , n7611 , n7612 );
not ( n7614 , n32 );
and ( n7615 , n7614 , n7604 );
nor ( n7616 , n7613 , n7615 );
nand ( n7617 , n7610 , n7616 );
nand ( n7618 , n35 , n7617 );
nand ( n7619 , n7606 , n7618 );
not ( n7620 , n7619 );
or ( n7621 , n7597 , n7620 );
nand ( n7622 , n7621 , n7377 );
nand ( n7623 , n724 , n7622 );
nand ( n7624 , n7595 , n7596 , n7623 );
and ( n7625 , n7624 , n2879 , n7519 );
not ( n7626 , n24 );
not ( n7627 , n534 );
not ( n7628 , n7528 );
or ( n7629 , n7627 , n7628 );
nand ( n7630 , n7629 , n7478 );
nand ( n7631 , n554 , n7630 );
nand ( n7632 , n554 , n7363 );
not ( n7633 , n35 );
nand ( n7634 , n7484 , n7578 );
not ( n7635 , n7634 );
not ( n7636 , n7536 );
or ( n7637 , n7635 , n7636 );
not ( n7638 , n32 );
and ( n7639 , n7638 , n7630 );
and ( n7640 , n927 , n7346 );
nor ( n7641 , n7639 , n7640 );
nand ( n7642 , n7637 , n7641 );
nand ( n7643 , n7633 , n7642 );
nand ( n7644 , n7631 , n7632 , n7643 );
not ( n7645 , n7644 );
or ( n7646 , n7626 , n7645 );
nand ( n7647 , n7646 , n7377 );
and ( n7648 , n7647 , n7380 , n3413 );
nor ( n7649 , n7625 , n7648 );
and ( n7650 , n7419 , n7518 , n7565 , n7649 );
not ( n7651 , n2458 );
nor ( n7652 , n7651 , n7416 );
and ( n7653 , n7380 , n7652 );
not ( n7654 , n1482 );
nand ( n7655 , n34 , n7426 );
not ( n7656 , n7473 );
nand ( n7657 , n7452 , n7655 , n7656 );
not ( n7658 , n7657 );
not ( n7659 , n7658 );
not ( n7660 , n7659 );
or ( n7661 , n7654 , n7660 );
nand ( n7662 , n7598 , n7428 );
nand ( n7663 , n7661 , n7662 );
or ( n7664 , n7363 , n7663 );
nand ( n7665 , n7664 , n7440 );
not ( n7666 , n35 );
not ( n7667 , n7486 );
nand ( n7668 , n382 , n7657 );
nand ( n7669 , n7496 , n7668 );
not ( n7670 , n7669 );
or ( n7671 , n7667 , n7670 );
not ( n7672 , n32 );
and ( n7673 , n7672 , n7663 );
nor ( n7674 , n895 , n7429 );
nor ( n7675 , n7673 , n7674 );
nand ( n7676 , n7671 , n7675 );
nand ( n7677 , n7666 , n7676 );
nand ( n7678 , n7665 , n7677 );
not ( n7679 , n7678 );
not ( n7680 , n24 );
or ( n7681 , n7679 , n7680 );
nand ( n7682 , n7681 , n7377 );
and ( n7683 , n3090 , n7380 , n3082 , n7682 );
not ( n7684 , n24 );
not ( n7685 , n7522 );
nand ( n7686 , n7526 , n7475 );
nor ( n7687 , n7530 , n7495 );
nand ( n7688 , n7686 , n7687 , n7497 );
nand ( n7689 , n7685 , n7688 );
and ( n7690 , n7494 , n7541 , n7497 , n7689 );
or ( n7691 , n7684 , n7690 );
nand ( n7692 , n7691 , n7377 );
and ( n7693 , n7519 , n2802 , n7692 );
nor ( n7694 , n7653 , n7683 , n7693 );
nor ( n7695 , n42 , n963 );
and ( n7696 , n7695 , n7396 );
and ( n7697 , n1919 , n7415 );
nor ( n7698 , n7696 , n7697 );
not ( n7699 , n2977 );
not ( n7700 , n7396 );
or ( n7701 , n7699 , n7700 );
nand ( n7702 , n7701 , n7556 );
nand ( n7703 , n908 , n7702 );
nand ( n7704 , n7698 , n7703 );
nand ( n7705 , n7380 , n7704 );
nor ( n7706 , n6723 , n7379 );
not ( n7707 , n24 );
not ( n7708 , n34 );
not ( n7709 , n7426 );
or ( n7710 , n7708 , n7709 );
nand ( n7711 , n7710 , n7527 );
and ( n7712 , n7526 , n7711 );
nor ( n7713 , n7712 , n7530 );
or ( n7714 , n7522 , n7713 );
and ( n7715 , n236 , n7711 );
nand ( n7716 , n7489 , n7535 );
nor ( n7717 , n7715 , n7716 );
buf ( n7718 , n7717 );
nand ( n7719 , n7714 , n7540 , n7718 );
not ( n7720 , n7719 );
or ( n7721 , n7707 , n7720 );
nand ( n7722 , n7721 , n7377 );
and ( n7723 , n590 , n7722 );
nor ( n7724 , n7723 , n7557 );
not ( n7725 , n24 );
not ( n7726 , n7522 );
nand ( n7727 , n7526 , n7659 );
nand ( n7728 , n7727 , n7687 , n7668 );
and ( n7729 , n7726 , n7728 );
nand ( n7730 , n7494 , n7541 );
not ( n7731 , n7668 );
nor ( n7732 , n7729 , n7730 , n7731 );
or ( n7733 , n7725 , n7732 );
nand ( n7734 , n7733 , n7377 );
nand ( n7735 , n520 , n7734 );
not ( n7736 , n24 );
not ( n7737 , n256 );
not ( n7738 , n7600 );
not ( n7739 , n7658 );
not ( n7740 , n7739 );
or ( n7741 , n7738 , n7740 );
not ( n7742 , n7427 );
nand ( n7743 , n1481 , n7742 );
nand ( n7744 , n7741 , n7743 );
not ( n7745 , n7744 );
nand ( n7746 , n7433 , n7745 );
not ( n7747 , n7746 );
or ( n7748 , n7737 , n7747 );
not ( n7749 , n7607 );
not ( n7750 , n7669 );
or ( n7751 , n7749 , n7750 );
not ( n7752 , n32 );
nand ( n7753 , n7752 , n7744 );
nand ( n7754 , n466 , n7430 );
nand ( n7755 , n7751 , n7753 , n7754 );
nand ( n7756 , n35 , n7755 );
nand ( n7757 , n7748 , n7756 );
not ( n7758 , n7757 );
or ( n7759 , n7736 , n7758 );
nand ( n7760 , n7759 , n7377 );
and ( n7761 , n724 , n7760 );
not ( n7762 , n24 );
not ( n7763 , n7598 );
not ( n7764 , n7711 );
or ( n7765 , n7763 , n7764 );
nand ( n7766 , n7765 , n7743 );
nand ( n7767 , n256 , n7766 );
not ( n7768 , n7579 );
or ( n7769 , n7768 , n7717 );
not ( n7770 , n32 );
nand ( n7771 , n7770 , n7766 );
nand ( n7772 , n216 , n7430 );
nand ( n7773 , n7769 , n7771 , n7772 );
nand ( n7774 , n35 , n7773 );
nand ( n7775 , n7767 , n7573 , n7774 );
not ( n7776 , n7775 );
or ( n7777 , n7762 , n7776 );
nand ( n7778 , n7777 , n7377 );
and ( n7779 , n96 , n7778 );
nor ( n7780 , n7761 , n7779 );
nand ( n7781 , n7724 , n7735 , n7780 );
not ( n7782 , n7781 );
buf ( n7783 , n7782 );
not ( n7784 , n7783 );
and ( n7785 , n7706 , n20 , n7784 );
nand ( n7786 , n16 , n2189 , n7415 );
nand ( n7787 , n2303 , n782 , n7396 );
nand ( n7788 , n2189 , n7702 );
nand ( n7789 , n7786 , n7787 , n7788 );
and ( n7790 , n7380 , n7789 );
nor ( n7791 , n7785 , n7790 );
not ( n7792 , n2 );
nand ( n7793 , n7792 , n1851 );
not ( n7794 , n7793 );
not ( n7795 , n7554 );
or ( n7796 , n7550 , n7795 );
nand ( n7797 , n7796 , n14 );
not ( n7798 , n7412 );
or ( n7799 , n7798 , n7403 );
not ( n7800 , n14 );
nand ( n7801 , n7799 , n7800 );
nand ( n7802 , n7797 , n2303 , n7801 );
not ( n7803 , n13 );
nor ( n7804 , n7803 , n1575 );
not ( n7805 , n7804 );
nand ( n7806 , n24 , n43 );
not ( n7807 , n7806 );
nand ( n7808 , n7807 , n7389 );
not ( n7809 , n43 );
nand ( n7810 , n5061 , n149 );
not ( n7811 , n7810 );
nand ( n7812 , n7809 , n7811 , n7373 );
nand ( n7813 , n7368 , n7808 , n7812 );
not ( n7814 , n7813 );
or ( n7815 , n1873 , n7814 );
not ( n7816 , n16 );
nand ( n7817 , n7816 , n7557 );
nand ( n7818 , n7815 , n7817 );
not ( n7819 , n7818 );
not ( n7820 , n24 );
and ( n7821 , n43 , n7820 , n4323 );
not ( n7822 , n7821 );
nor ( n7823 , n632 , n7822 );
not ( n7824 , n1482 );
not ( n7825 , n7455 );
not ( n7826 , n7354 );
not ( n7827 , n7826 );
or ( n7828 , n7825 , n7827 );
not ( n7829 , n7337 );
nor ( n7830 , n7444 , n7829 );
not ( n7831 , n7359 );
nor ( n7832 , n7830 , n7831 );
nand ( n7833 , n7828 , n7832 );
nand ( n7834 , n34 , n7833 );
not ( n7835 , n36 );
not ( n7836 , n7360 );
or ( n7837 , n7835 , n7836 );
not ( n7838 , n36 );
not ( n7839 , n7833 );
and ( n7840 , n7838 , n7839 );
nor ( n7841 , n7840 , n34 );
nand ( n7842 , n7837 , n7841 );
nand ( n7843 , n7834 , n7842 );
not ( n7844 , n7843 );
or ( n7845 , n7824 , n7844 );
not ( n7846 , n7598 );
not ( n7847 , n7833 );
or ( n7848 , n7846 , n7847 );
nand ( n7849 , n7845 , n7848 );
nand ( n7850 , n7440 , n7849 );
not ( n7851 , n26 );
and ( n7852 , n234 , n7386 );
nand ( n7853 , n7851 , n7852 );
nand ( n7854 , n7352 , n7853 );
nand ( n7855 , n7440 , n7854 );
not ( n7856 , n35 );
nand ( n7857 , n232 , n7852 );
nand ( n7858 , n7484 , n7857 );
not ( n7859 , n7858 );
not ( n7860 , n236 );
not ( n7861 , n7843 );
or ( n7862 , n7860 , n7861 );
and ( n7863 , n7534 , n7852 );
not ( n7864 , n7489 );
nor ( n7865 , n7863 , n7864 );
nand ( n7866 , n7862 , n7865 );
not ( n7867 , n7866 );
or ( n7868 , n7859 , n7867 );
not ( n7869 , n32 );
and ( n7870 , n7869 , n7849 );
not ( n7871 , n7847 );
not ( n7872 , n7871 );
nor ( n7873 , n607 , n7872 );
nor ( n7874 , n7870 , n7873 );
nand ( n7875 , n7868 , n7874 );
nand ( n7876 , n7856 , n7875 );
nand ( n7877 , n7850 , n7855 , n7876 );
and ( n7878 , n7823 , n7877 );
nor ( n7879 , n521 , n7822 );
not ( n7880 , n7854 );
not ( n7881 , n7880 );
not ( n7882 , n1482 );
not ( n7883 , n34 );
not ( n7884 , n7833 );
or ( n7885 , n7883 , n7884 );
not ( n7886 , n34 );
not ( n7887 , n7422 );
nand ( n7888 , n7886 , n393 , n7887 );
and ( n7889 , n7463 , n7888 );
nand ( n7890 , n7885 , n7889 );
not ( n7891 , n7890 );
or ( n7892 , n7882 , n7891 );
nand ( n7893 , n7892 , n7848 );
not ( n7894 , n7893 );
not ( n7895 , n7894 );
or ( n7896 , n7881 , n7895 );
nand ( n7897 , n7896 , n7440 );
not ( n7898 , n35 );
nand ( n7899 , n37 , n7852 );
and ( n7900 , n7484 , n7899 );
not ( n7901 , n382 );
not ( n7902 , n7890 );
or ( n7903 , n7901 , n7902 );
nand ( n7904 , n7493 , n7852 );
and ( n7905 , n7489 , n7904 );
nand ( n7906 , n7903 , n7905 );
not ( n7907 , n7906 );
or ( n7908 , n7900 , n7907 );
or ( n7909 , n32 , n7894 );
nand ( n7910 , n531 , n7871 );
nand ( n7911 , n7908 , n7909 , n7910 );
nand ( n7912 , n7898 , n7911 );
nand ( n7913 , n7897 , n7912 );
and ( n7914 , n7879 , n7913 );
nor ( n7915 , n7878 , n7914 );
nand ( n7916 , n7819 , n7915 );
not ( n7917 , n24 );
nor ( n7918 , n7917 , n22 );
not ( n7919 , n7918 );
or ( n7920 , n43 , n7919 );
nor ( n7921 , n7920 , n632 );
not ( n7922 , n7921 );
not ( n7923 , n7439 );
not ( n7924 , n1481 );
not ( n7925 , n7711 );
or ( n7926 , n7924 , n7925 );
nand ( n7927 , n7926 , n7662 );
nand ( n7928 , n7923 , n7927 );
not ( n7929 , n7634 );
nor ( n7930 , n7929 , n7717 );
not ( n7931 , n7927 );
or ( n7932 , n32 , n7931 );
not ( n7933 , n7429 );
nand ( n7934 , n927 , n7933 );
nand ( n7935 , n7932 , n7934 );
or ( n7936 , n7930 , n7935 );
not ( n7937 , n35 );
nand ( n7938 , n7936 , n7937 );
nand ( n7939 , n7928 , n7632 , n7938 );
not ( n7940 , n7939 );
or ( n7941 , n7922 , n7940 );
nor ( n7942 , n7920 , n521 );
nand ( n7943 , n7942 , n7678 );
nand ( n7944 , n7941 , n7943 );
nor ( n7945 , n7916 , n7944 );
or ( n7946 , n7805 , n7945 );
not ( n7947 , n20 );
not ( n7948 , n19 );
nand ( n7949 , n13 , n18 );
not ( n7950 , n7949 );
nand ( n7951 , n7948 , n7950 );
nor ( n7952 , n7947 , n7951 );
not ( n7953 , n7952 );
not ( n7954 , n3434 );
not ( n7955 , n7814 );
and ( n7956 , n7954 , n7955 );
not ( n7957 , n7596 );
nor ( n7958 , n7956 , n7957 );
nor ( n7959 , n295 , n7822 );
not ( n7960 , n7599 );
not ( n7961 , n7960 );
not ( n7962 , n7843 );
or ( n7963 , n7961 , n7962 );
not ( n7964 , n1481 );
or ( n7965 , n7964 , n7847 );
nand ( n7966 , n7963 , n7965 );
nand ( n7967 , n256 , n7966 );
nand ( n7968 , n256 , n7854 );
not ( n7969 , n32 );
nand ( n7970 , n7969 , n7966 );
not ( n7971 , n7970 );
not ( n7972 , n215 );
not ( n7973 , n7872 );
and ( n7974 , n7972 , n7973 );
nand ( n7975 , n7575 , n7857 );
and ( n7976 , n7975 , n7866 );
nor ( n7977 , n7974 , n7976 );
not ( n7978 , n7977 );
or ( n7979 , n7971 , n7978 );
nand ( n7980 , n7979 , n35 );
nand ( n7981 , n7967 , n7968 , n7980 );
and ( n7982 , n7959 , n7981 );
nor ( n7983 , n1316 , n7822 );
not ( n7984 , n7960 );
not ( n7985 , n7890 );
or ( n7986 , n7984 , n7985 );
nand ( n7987 , n7986 , n7965 );
or ( n7988 , n7854 , n7987 );
nand ( n7989 , n7988 , n256 );
not ( n7990 , n32 );
nand ( n7991 , n7990 , n7987 );
nand ( n7992 , n466 , n7871 );
nand ( n7993 , n7575 , n7899 );
nand ( n7994 , n7993 , n7906 );
and ( n7995 , n7991 , n7992 , n7994 );
not ( n7996 , n35 );
nor ( n7997 , n7995 , n7996 );
not ( n7998 , n7997 );
nand ( n7999 , n7989 , n7998 );
and ( n8000 , n7983 , n7999 );
nor ( n8001 , n7982 , n8000 );
nand ( n8002 , n7958 , n8001 );
nor ( n8003 , n7920 , n295 );
not ( n8004 , n8003 );
not ( n8005 , n7775 );
or ( n8006 , n8004 , n8005 );
nor ( n8007 , n7920 , n1316 );
nand ( n8008 , n8007 , n7757 );
nand ( n8009 , n8006 , n8008 );
nor ( n8010 , n8002 , n8009 );
or ( n8011 , n7953 , n8010 );
nand ( n8012 , n7946 , n8011 );
nand ( n8013 , n7802 , n8012 );
not ( n8014 , n7685 );
nand ( n8015 , n7526 , n7890 );
and ( n8016 , n8015 , n7531 , n7907 );
or ( n8017 , n8014 , n8016 );
and ( n8018 , n1382 , n7852 );
nor ( n8019 , n8018 , n7906 );
nand ( n8020 , n8017 , n8019 );
not ( n8021 , n8020 );
nand ( n8022 , n13 , n1582 );
nor ( n8023 , n8021 , n8022 );
not ( n8024 , n2306 );
and ( n8025 , n8023 , n7811 , n8024 );
not ( n8026 , n2937 );
not ( n8027 , n8022 );
nand ( n8028 , n8026 , n8027 , n3299 , n7811 );
not ( n8029 , n17 );
not ( n8030 , n7843 );
or ( n8031 , n7525 , n8030 );
nand ( n8032 , n8031 , n7531 );
and ( n8033 , n7685 , n8032 );
not ( n8034 , n7853 );
and ( n8035 , n32 , n8034 );
nor ( n8036 , n8033 , n8035 , n7866 );
nor ( n8037 , n8028 , n8029 , n8036 );
nor ( n8038 , n8025 , n8037 );
and ( n8039 , n7389 , n7918 , n149 );
nor ( n8040 , n8039 , n7367 );
or ( n8041 , n42 , n8040 );
or ( n8042 , n795 , n8041 );
not ( n8043 , n16 );
and ( n8044 , n8043 , n6725 );
and ( n8045 , n8044 , n7413 );
and ( n8046 , n3299 , n7795 );
nor ( n8047 , n8045 , n8046 );
nand ( n8048 , n8042 , n8047 );
nand ( n8049 , n8027 , n8048 );
not ( n8050 , n8041 );
nand ( n8051 , n8050 , n3185 , n3352 );
or ( n8052 , n1891 , n8041 );
nand ( n8053 , n8052 , n7551 );
nand ( n8054 , n3146 , n8053 );
nor ( n8055 , n972 , n8041 );
nand ( n8056 , n453 , n8055 );
not ( n8057 , n8055 );
nand ( n8058 , n8057 , n7596 );
nand ( n8059 , n629 , n8058 );
nand ( n8060 , n8051 , n8054 , n8056 , n8059 );
or ( n8061 , n42 , n7810 );
not ( n8062 , n8061 );
nand ( n8063 , n8062 , n2255 );
not ( n8064 , n7880 );
not ( n8065 , n7960 );
nand ( n8066 , n34 , n7361 );
nand ( n8067 , n7889 , n8066 );
not ( n8068 , n8067 );
or ( n8069 , n8065 , n8068 );
not ( n8070 , n34 );
not ( n8071 , n8070 );
not ( n8072 , n7833 );
or ( n8073 , n8071 , n8072 );
nand ( n8074 , n8073 , n8066 );
nand ( n8075 , n1482 , n8074 );
nand ( n8076 , n8069 , n8075 );
not ( n8077 , n8076 );
not ( n8078 , n8077 );
or ( n8079 , n8064 , n8078 );
nand ( n8080 , n8079 , n256 );
not ( n8081 , n32 );
nand ( n8082 , n8081 , n8076 );
not ( n8083 , n8082 );
not ( n8084 , n382 );
not ( n8085 , n8067 );
or ( n8086 , n8084 , n8085 );
nand ( n8087 , n8086 , n7905 );
and ( n8088 , n7993 , n8087 );
and ( n8089 , n466 , n8074 );
nor ( n8090 , n8088 , n8089 );
not ( n8091 , n8090 );
or ( n8092 , n8083 , n8091 );
nand ( n8093 , n8092 , n35 );
nand ( n8094 , n8080 , n8093 );
not ( n8095 , n8094 );
or ( n8096 , n8063 , n8095 );
nand ( n8097 , n8062 , n522 );
not ( n8098 , n7440 );
not ( n8099 , n1482 );
not ( n8100 , n8067 );
or ( n8101 , n8099 , n8100 );
nand ( n8102 , n7600 , n8074 );
nand ( n8103 , n8101 , n8102 );
not ( n8104 , n8103 );
nand ( n8105 , n8104 , n7880 );
not ( n8106 , n8105 );
or ( n8107 , n8098 , n8106 );
not ( n8108 , n35 );
not ( n8109 , n7900 );
nand ( n8110 , n8109 , n8087 );
nand ( n8111 , n531 , n8074 );
not ( n8112 , n32 );
nand ( n8113 , n8112 , n8103 );
nand ( n8114 , n8110 , n8111 , n8113 );
nand ( n8115 , n8108 , n8114 );
nand ( n8116 , n8107 , n8115 );
not ( n8117 , n8116 );
or ( n8118 , n8097 , n8117 );
not ( n8119 , n8067 );
or ( n8120 , n8119 , n7525 );
nand ( n8121 , n8120 , n7531 );
and ( n8122 , n7726 , n8121 );
nor ( n8123 , n8122 , n8035 , n8087 );
not ( n8124 , n8123 );
not ( n8125 , n6283 );
and ( n8126 , n8124 , n8062 , n8125 );
or ( n8127 , n6283 , n8041 );
or ( n8128 , n20 , n8047 );
nand ( n8129 , n8127 , n8128 );
nor ( n8130 , n8126 , n8129 );
nand ( n8131 , n8096 , n8118 , n8130 );
or ( n8132 , n8060 , n8131 );
not ( n8133 , n7920 );
and ( n8134 , n8133 , n7543 );
not ( n8135 , n7526 );
nand ( n8136 , n8066 , n7842 );
not ( n8137 , n8136 );
or ( n8138 , n8135 , n8137 );
nand ( n8139 , n8138 , n7531 );
nand ( n8140 , n7685 , n8139 );
not ( n8141 , n8035 );
not ( n8142 , n236 );
not ( n8143 , n8136 );
or ( n8144 , n8142 , n8143 );
nand ( n8145 , n8144 , n7865 );
not ( n8146 , n8145 );
and ( n8147 , n8140 , n8141 , n8146 );
nor ( n8148 , n7822 , n8147 );
nor ( n8149 , n8134 , n8148 , n7813 );
or ( n8150 , n3182 , n8149 );
nor ( n8151 , n571 , n8061 );
not ( n8152 , n8151 );
not ( n8153 , n8074 );
not ( n8154 , n8153 );
and ( n8155 , n8154 , n25 );
nor ( n8156 , n8155 , n7854 );
or ( n8157 , n8152 , n8156 );
nand ( n8158 , n8150 , n8157 );
not ( n8159 , n2190 );
and ( n8160 , n8159 , n7802 );
not ( n8161 , n8160 );
and ( n8162 , n7942 , n7510 );
and ( n8163 , n7879 , n8116 );
nor ( n8164 , n8162 , n8163 );
not ( n8165 , n7645 );
nand ( n8166 , n8165 , n7921 );
not ( n8167 , n32 );
not ( n8168 , n1482 );
not ( n8169 , n8136 );
or ( n8170 , n8168 , n8169 );
nand ( n8171 , n8170 , n8102 );
and ( n8172 , n8167 , n8171 );
not ( n8173 , n7858 );
not ( n8174 , n8145 );
or ( n8175 , n8173 , n8174 );
not ( n8176 , n8153 );
nand ( n8177 , n927 , n8176 );
nand ( n8178 , n8175 , n8177 );
or ( n8179 , n8172 , n8178 );
not ( n8180 , n35 );
nand ( n8181 , n8179 , n8180 );
nand ( n8182 , n7440 , n8171 );
nand ( n8183 , n8181 , n7855 , n8182 );
nand ( n8184 , n7823 , n8183 );
nand ( n8185 , n8164 , n7819 , n8166 , n8184 );
not ( n8186 , n8185 );
or ( n8187 , n8161 , n8186 );
not ( n8188 , n2408 );
or ( n8189 , n7822 , n8156 );
or ( n8190 , n7920 , n7364 );
nand ( n8191 , n8189 , n8190 , n7814 );
nand ( n8192 , n8188 , n8191 , n2191 );
nand ( n8193 , n8187 , n8192 );
nor ( n8194 , n8158 , n8193 );
or ( n8195 , n7920 , n7690 );
or ( n8196 , n7822 , n8123 );
nand ( n8197 , n8195 , n8196 , n7814 );
and ( n8198 , n2418 , n8197 );
nor ( n8199 , n2446 , n3493 , n8061 );
not ( n8200 , n8147 );
and ( n8201 , n8199 , n8200 );
nor ( n8202 , n8198 , n8201 );
nand ( n8203 , n8062 , n1571 );
not ( n8204 , n8183 );
nor ( n8205 , n8203 , n8204 );
and ( n8206 , n8007 , n7619 );
and ( n8207 , n7983 , n8094 );
nor ( n8208 , n8206 , n8207 );
not ( n8209 , n7960 );
not ( n8210 , n8136 );
or ( n8211 , n8209 , n8210 );
nand ( n8212 , n8211 , n8075 );
nand ( n8213 , n256 , n8212 );
not ( n8214 , n32 );
and ( n8215 , n8214 , n8212 );
not ( n8216 , n7975 );
not ( n8217 , n8145 );
or ( n8218 , n8216 , n8217 );
nand ( n8219 , n216 , n8074 );
nand ( n8220 , n8218 , n8219 );
or ( n8221 , n8215 , n8220 );
nand ( n8222 , n8221 , n35 );
nand ( n8223 , n8213 , n7968 , n8222 );
and ( n8224 , n7959 , n8223 );
and ( n8225 , n8003 , n7591 );
nor ( n8226 , n8224 , n8225 );
and ( n8227 , n8208 , n7958 , n8226 );
nand ( n8228 , n453 , n7802 );
or ( n8229 , n8227 , n8228 );
nand ( n8230 , n8062 , n842 );
not ( n8231 , n8223 );
or ( n8232 , n8230 , n8231 );
nand ( n8233 , n8229 , n8232 );
nor ( n8234 , n8205 , n8233 );
nand ( n8235 , n8194 , n8202 , n8234 );
or ( n8236 , n8132 , n8235 );
nand ( n8237 , n8236 , n7950 );
and ( n8238 , n8013 , n8038 , n8049 , n8237 );
and ( n8239 , n8133 , n7719 );
nor ( n8240 , n7822 , n8036 );
nor ( n8241 , n8239 , n8240 , n7813 );
or ( n8242 , n8241 , n8022 , n3309 );
not ( n8243 , n7981 );
nand ( n8244 , n7952 , n8062 );
or ( n8245 , n8243 , n295 , n8244 );
nand ( n8246 , n8242 , n8245 );
not ( n8247 , n8246 );
and ( n8248 , n8053 , n8027 , n3299 );
nor ( n8249 , n234 , n7847 );
nor ( n8250 , n7854 , n8249 );
buf ( n8251 , n3436 );
nand ( n8252 , n7804 , n8062 );
nor ( n8253 , n8250 , n8251 , n8252 );
nor ( n8254 , n8248 , n8253 );
and ( n8255 , n7804 , n8058 );
and ( n8256 , n7952 , n8055 );
nor ( n8257 , n8255 , n8256 );
nand ( n8258 , n8247 , n8254 , n8257 );
not ( n8259 , n7999 );
or ( n8260 , n8259 , n1316 , n8244 );
not ( n8261 , n7913 );
or ( n8262 , n8261 , n521 , n8252 );
nand ( n8263 , n8260 , n8262 );
and ( n8264 , n8133 , n7434 );
nor ( n8265 , n7822 , n8250 );
nor ( n8266 , n8264 , n8265 , n7813 );
or ( n8267 , n8266 , n2408 , n7805 );
or ( n8268 , n8041 , n1873 , n7805 );
nand ( n8269 , n8267 , n8268 );
and ( n8270 , n7821 , n8020 );
or ( n8271 , n7920 , n7732 );
nand ( n8272 , n8271 , n7814 );
nor ( n8273 , n8270 , n8272 );
or ( n8274 , n8273 , n8022 , n2450 );
not ( n8275 , n7877 );
or ( n8276 , n8275 , n632 , n8252 );
nand ( n8277 , n8274 , n8276 );
nor ( n8278 , n8258 , n8263 , n8269 , n8277 );
and ( n8279 , n908 , n7802 );
buf ( n8280 , n1105 );
not ( n8281 , n8280 );
and ( n8282 , n8281 , n7663 );
not ( n8283 , n7677 );
not ( n8284 , n1306 );
not ( n8285 , n7430 );
or ( n8286 , n8284 , n8285 );
nand ( n8287 , n8286 , n7531 );
nor ( n8288 , n8282 , n8283 , n8287 );
not ( n8289 , n32 );
and ( n8290 , n8289 , n7678 );
not ( n8291 , n1651 );
not ( n8292 , n8291 );
not ( n8293 , n8292 );
not ( n8294 , n8293 );
not ( n8295 , n8294 );
and ( n8296 , n8295 , n7659 );
nor ( n8297 , n8290 , n8296 );
nand ( n8298 , n8288 , n8297 );
and ( n8299 , n7942 , n8298 );
nor ( n8300 , n8299 , n7818 );
and ( n8301 , n8281 , n7927 );
nor ( n8302 , n8301 , n8287 );
not ( n8303 , n32 );
and ( n8304 , n8303 , n7939 );
and ( n8305 , n8293 , n7711 );
nor ( n8306 , n8304 , n8305 );
nand ( n8307 , n8302 , n7938 , n8306 );
nand ( n8308 , n7921 , n8307 );
not ( n8309 , n32 );
not ( n8310 , n8275 );
and ( n8311 , n8309 , n8310 );
not ( n8312 , n7876 );
nor ( n8313 , n8311 , n8312 );
not ( n8314 , n7872 );
and ( n8315 , n1306 , n8314 );
nor ( n8316 , n8315 , n7530 );
not ( n8317 , n8280 );
not ( n8318 , n8317 );
not ( n8319 , n8318 );
and ( n8320 , n8319 , n7849 );
not ( n8321 , n8294 );
not ( n8322 , n8030 );
and ( n8323 , n8321 , n8322 );
nor ( n8324 , n8320 , n8323 );
nand ( n8325 , n8313 , n8316 , n8324 );
and ( n8326 , n7823 , n8325 );
or ( n8327 , n8318 , n7894 );
nand ( n8328 , n8327 , n8316 );
not ( n8329 , n7912 );
nor ( n8330 , n8328 , n8329 );
not ( n8331 , n32 );
and ( n8332 , n8331 , n7913 );
and ( n8333 , n8321 , n7890 );
nor ( n8334 , n8332 , n8333 );
nand ( n8335 , n8330 , n8334 );
and ( n8336 , n7879 , n8335 );
nor ( n8337 , n8326 , n8336 );
nand ( n8338 , n8300 , n8308 , n8337 );
and ( n8339 , n8279 , n8338 );
nor ( n8340 , n912 , n8061 );
and ( n8341 , n8325 , n590 , n8340 );
nor ( n8342 , n8339 , n8341 );
or ( n8343 , n8280 , n7745 );
and ( n8344 , n8291 , n7430 );
nor ( n8345 , n8344 , n7530 );
nand ( n8346 , n8343 , n8345 );
not ( n8347 , n7756 );
nor ( n8348 , n8346 , n8347 );
not ( n8349 , n1306 );
not ( n8350 , n8349 );
not ( n8351 , n8350 );
not ( n8352 , n8351 );
nand ( n8353 , n8352 , n7659 );
not ( n8354 , n32 );
nand ( n8355 , n8354 , n7757 );
nand ( n8356 , n8348 , n8353 , n8355 );
and ( n8357 , n8007 , n8356 );
not ( n8358 , n7958 );
nor ( n8359 , n8357 , n8358 );
and ( n8360 , n8319 , n7966 );
and ( n8361 , n8352 , n8322 );
nor ( n8362 , n8360 , n8361 );
or ( n8363 , n8292 , n7872 );
nand ( n8364 , n8363 , n7531 );
or ( n8365 , n32 , n8243 );
nand ( n8366 , n8365 , n7980 );
nor ( n8367 , n8364 , n8366 );
nand ( n8368 , n8362 , n8367 );
and ( n8369 , n7959 , n8368 );
not ( n8370 , n8280 );
and ( n8371 , n8370 , n7987 );
nor ( n8372 , n8371 , n7997 , n8364 );
not ( n8373 , n32 );
and ( n8374 , n8373 , n7999 );
and ( n8375 , n8352 , n7890 );
nor ( n8376 , n8374 , n8375 );
nand ( n8377 , n8372 , n8376 );
and ( n8378 , n7983 , n8377 );
nor ( n8379 , n8369 , n8378 );
and ( n8380 , n8281 , n7766 );
not ( n8381 , n8345 );
nor ( n8382 , n8380 , n8381 );
not ( n8383 , n8351 );
not ( n8384 , n7711 );
not ( n8385 , n8384 );
and ( n8386 , n8383 , n8385 );
not ( n8387 , n32 );
and ( n8388 , n8387 , n7775 );
nor ( n8389 , n8386 , n8388 );
nand ( n8390 , n8382 , n7774 , n8389 );
nand ( n8391 , n8003 , n8390 );
and ( n8392 , n8359 , n8379 , n8391 );
nor ( n8393 , n8392 , n2439 );
nand ( n8394 , n7802 , n8393 );
not ( n8395 , n7475 );
or ( n8396 , n8294 , n8395 );
and ( n8397 , n8281 , n7479 );
nor ( n8398 , n8349 , n7502 );
nor ( n8399 , n8397 , n8398 , n7530 );
not ( n8400 , n32 );
and ( n8401 , n8400 , n7510 );
not ( n8402 , n7509 );
nor ( n8403 , n8401 , n8402 );
nand ( n8404 , n8396 , n8399 , n8403 );
and ( n8405 , n7942 , n8404 );
and ( n8406 , n8317 , n7630 );
nand ( n8407 , n8293 , n7528 );
not ( n8408 , n32 );
nand ( n8409 , n8408 , n7644 );
nand ( n8410 , n7643 , n8407 , n8409 );
nor ( n8411 , n8406 , n8410 );
not ( n8412 , n8398 );
nand ( n8413 , n8411 , n7531 , n8412 );
and ( n8414 , n7921 , n8413 );
nor ( n8415 , n8405 , n8414 );
nand ( n8416 , n32 , n8067 );
or ( n8417 , n1054 , n8416 );
not ( n8418 , n32 );
not ( n8419 , n8117 );
and ( n8420 , n8418 , n8419 );
not ( n8421 , n8115 );
nor ( n8422 , n8420 , n8421 );
and ( n8423 , n8317 , n8103 );
not ( n8424 , n8154 );
nor ( n8425 , n8351 , n8424 );
nor ( n8426 , n8423 , n7530 , n8425 );
nand ( n8427 , n8417 , n8422 , n8426 );
and ( n8428 , n7879 , n8427 );
not ( n8429 , n7823 );
and ( n8430 , n8321 , n8136 );
nor ( n8431 , n8430 , n7530 );
and ( n8432 , n8319 , n8171 );
nor ( n8433 , n8432 , n8425 );
not ( n8434 , n32 );
nand ( n8435 , n8434 , n8183 );
nand ( n8436 , n8431 , n8433 , n8181 , n8435 );
not ( n8437 , n8436 );
or ( n8438 , n8429 , n8437 );
nand ( n8439 , n8438 , n7819 );
nor ( n8440 , n8428 , n8439 );
nand ( n8441 , n8415 , n8440 );
nand ( n8442 , n8160 , n8441 );
nand ( n8443 , n8342 , n8394 , n8442 );
not ( n8444 , n8228 );
not ( n8445 , n8319 );
or ( n8446 , n8445 , n8077 );
nand ( n8447 , n8293 , n8154 );
not ( n8448 , n8447 );
or ( n8449 , n1442 , n8416 );
nand ( n8450 , n8449 , n7531 );
nor ( n8451 , n8448 , n8450 );
not ( n8452 , n32 );
and ( n8453 , n8452 , n8094 );
not ( n8454 , n8093 );
nor ( n8455 , n8453 , n8454 );
nand ( n8456 , n8446 , n8451 , n8455 );
and ( n8457 , n7983 , n8456 );
nor ( n8458 , n8292 , n7502 );
not ( n8459 , n8458 );
nand ( n8460 , n8317 , n7571 );
not ( n8461 , n7590 );
not ( n8462 , n32 );
not ( n8463 , n8462 );
not ( n8464 , n7591 );
or ( n8465 , n8463 , n8464 );
nand ( n8466 , n8350 , n7528 );
nand ( n8467 , n8465 , n8466 );
nor ( n8468 , n8461 , n8467 );
nand ( n8469 , n7531 , n8459 , n8460 , n8468 );
and ( n8470 , n8003 , n8469 );
nor ( n8471 , n8457 , n8470 );
not ( n8472 , n8280 );
and ( n8473 , n8472 , n7604 );
nor ( n8474 , n8473 , n8458 , n7530 );
nand ( n8475 , n8352 , n7475 );
not ( n8476 , n32 );
nand ( n8477 , n8476 , n7619 );
nand ( n8478 , n8474 , n8475 , n7618 , n8477 );
nand ( n8479 , n8007 , n8478 );
and ( n8480 , n8352 , n8136 );
nor ( n8481 , n8480 , n7530 );
not ( n8482 , n8319 );
not ( n8483 , n8212 );
or ( n8484 , n8482 , n8483 );
nand ( n8485 , n8484 , n8447 );
not ( n8486 , n32 );
not ( n8487 , n8486 );
not ( n8488 , n8223 );
or ( n8489 , n8487 , n8488 );
nand ( n8490 , n8489 , n8222 );
nor ( n8491 , n8485 , n8490 );
nand ( n8492 , n8481 , n8491 );
nand ( n8493 , n7959 , n8492 );
nand ( n8494 , n8471 , n8479 , n7958 , n8493 );
and ( n8495 , n8444 , n8494 );
not ( n8496 , n8456 );
nor ( n8497 , n8063 , n8496 );
nor ( n8498 , n8495 , n8497 );
not ( n8499 , n2434 );
nor ( n8500 , n8499 , n8061 );
and ( n8501 , n8368 , n96 , n8500 );
and ( n8502 , n8335 , n520 , n8340 );
nor ( n8503 , n8501 , n8502 );
or ( n8504 , n32 , n8156 );
or ( n8505 , n7525 , n8424 );
nand ( n8506 , n8504 , n8505 , n7531 );
and ( n8507 , n7821 , n8506 );
or ( n8508 , n32 , n7364 );
or ( n8509 , n7525 , n7502 );
nand ( n8510 , n8508 , n8509 , n7531 );
not ( n8511 , n8510 );
or ( n8512 , n7920 , n8511 );
nand ( n8513 , n8512 , n7814 );
nor ( n8514 , n8507 , n8513 );
or ( n8515 , n8514 , n2192 , n2408 );
nand ( n8516 , n8515 , n8054 );
and ( n8517 , n8377 , n724 , n8500 );
not ( n8518 , n7811 );
nor ( n8519 , n8032 , n7866 );
nor ( n8520 , n8518 , n2391 , n8519 , n2396 );
nor ( n8521 , n8517 , n8520 );
or ( n8522 , n8121 , n8087 );
nand ( n8523 , n8062 , n8125 , n8522 );
nand ( n8524 , n8059 , n8523 );
nand ( n8525 , n7713 , n7718 );
nand ( n8526 , n8133 , n8525 );
or ( n8527 , n7822 , n8519 );
and ( n8528 , n8526 , n7814 , n8527 );
or ( n8529 , n2431 , n8528 );
not ( n8530 , n2409 );
not ( n8531 , n32 );
and ( n8532 , n8531 , n7434 );
or ( n8533 , n7525 , n8285 );
nand ( n8534 , n8533 , n7531 );
nor ( n8535 , n8532 , n8534 );
or ( n8536 , n8535 , n7920 );
or ( n8537 , n32 , n8250 );
or ( n8538 , n7525 , n7847 );
nand ( n8539 , n8537 , n8538 , n7531 );
nand ( n8540 , n7821 , n8539 );
nand ( n8541 , n8536 , n7814 , n8540 );
not ( n8542 , n8541 );
or ( n8543 , n8530 , n8542 );
nand ( n8544 , n8529 , n8543 );
nor ( n8545 , n8524 , n8544 );
and ( n8546 , n7821 , n8522 );
not ( n8547 , n7688 );
or ( n8548 , n7920 , n8547 );
nand ( n8549 , n8548 , n7814 );
nor ( n8550 , n8546 , n8549 );
not ( n8551 , n8550 );
and ( n8552 , n2418 , n8551 );
not ( n8553 , n8139 );
nand ( n8554 , n8553 , n8146 );
and ( n8555 , n8199 , n8554 );
nor ( n8556 , n8552 , n8555 , n8129 );
and ( n8557 , n908 , n8058 );
or ( n8558 , n7822 , n8016 );
not ( n8559 , n7728 );
or ( n8560 , n7920 , n8559 );
nand ( n8561 , n8558 , n8560 , n7814 );
and ( n8562 , n3221 , n8561 );
and ( n8563 , n20 , n8048 );
and ( n8564 , n644 , n8055 );
nor ( n8565 , n8563 , n8564 );
not ( n8566 , n8565 );
nand ( n8567 , n20 , n2123 );
or ( n8568 , n8016 , n8061 , n8567 );
or ( n8569 , n8041 , n912 , n1873 );
nand ( n8570 , n8568 , n8569 );
nor ( n8571 , n8566 , n8570 );
not ( n8572 , n1960 );
and ( n8573 , n8539 , n8572 , n8340 );
and ( n8574 , n2392 , n8053 );
nor ( n8575 , n8573 , n8574 );
nand ( n8576 , n8571 , n8575 , n8051 , n8056 );
nor ( n8577 , n8557 , n8562 , n8576 );
nand ( n8578 , n8521 , n8545 , n8556 , n8577 );
nor ( n8579 , n8516 , n8578 );
not ( n8580 , n8097 );
and ( n8581 , n8580 , n8427 );
or ( n8582 , n7920 , n7538 );
nand ( n8583 , n7821 , n8554 );
nand ( n8584 , n8582 , n7814 , n8583 );
and ( n8585 , n2447 , n8584 );
nor ( n8586 , n8581 , n8585 );
not ( n8587 , n8492 );
not ( n8588 , n8587 );
not ( n8589 , n8230 );
and ( n8590 , n8588 , n8589 );
not ( n8591 , n8151 );
not ( n8592 , n8506 );
or ( n8593 , n8591 , n8592 );
not ( n8594 , n8436 );
or ( n8595 , n8203 , n8594 );
nand ( n8596 , n8593 , n8595 );
nor ( n8597 , n8590 , n8596 );
and ( n8598 , n8503 , n8579 , n8586 , n8597 );
nand ( n8599 , n8498 , n8598 );
or ( n8600 , n8443 , n8599 );
not ( n8601 , n13 );
nor ( n8602 , n8601 , n18 );
nand ( n8603 , n8600 , n8602 );
nand ( n8604 , n8238 , n8278 , n8603 );
nand ( n8605 , n7794 , n8604 );
and ( n8606 , n7694 , n7705 , n7791 , n8605 );
not ( n8607 , n993 );
nor ( n8608 , n3471 , n2791 );
not ( n8609 , n7806 );
not ( n8610 , n24 );
not ( n8611 , n8525 );
or ( n8612 , n8610 , n8611 );
nand ( n8613 , n8612 , n7377 );
not ( n8614 , n8613 );
or ( n8615 , n8609 , n8614 );
not ( n8616 , n4312 );
not ( n8617 , n8616 );
not ( n8618 , n8617 );
not ( n8619 , n8618 );
not ( n8620 , n8619 );
buf ( n8621 , n8620 );
not ( n8622 , n8621 );
or ( n8623 , n7806 , n8622 );
nand ( n8624 , n24 , n31 );
nand ( n8625 , n8624 , n7808 );
not ( n8626 , n8625 );
nand ( n8627 , n8623 , n8626 );
not ( n8628 , n8627 );
nand ( n8629 , n8615 , n8628 );
and ( n8630 , n8608 , n8629 );
nor ( n8631 , n2384 , n3471 );
not ( n8632 , n8631 );
nor ( n8633 , n16 , n1404 );
not ( n8634 , n8633 );
and ( n8635 , n8632 , n8634 );
nor ( n8636 , n8635 , n7416 );
not ( n8637 , n7563 );
not ( n8638 , n7789 );
and ( n8639 , n8637 , n8638 );
nor ( n8640 , n8639 , n18 );
nor ( n8641 , n8630 , n8636 , n8640 );
not ( n8642 , n24 );
not ( n8643 , n8619 );
or ( n8644 , n7809 , n8642 , n8643 );
not ( n8645 , n8644 );
and ( n8646 , n24 , n8404 );
nor ( n8647 , n8646 , n7376 );
or ( n8648 , n8645 , n8647 );
nand ( n8649 , n8648 , n8626 );
and ( n8650 , n8649 , n3082 , n8633 );
not ( n8651 , n18 );
and ( n8652 , n8651 , n7704 );
nor ( n8653 , n8650 , n8652 );
not ( n8654 , n18 );
not ( n8655 , n24 );
not ( n8656 , n8307 );
or ( n8657 , n8655 , n8656 );
nand ( n8658 , n8657 , n7377 );
and ( n8659 , n8658 , n8644 );
nor ( n8660 , n8659 , n8625 );
nor ( n8661 , n8660 , n913 );
nand ( n8662 , n42 , n8654 , n8661 );
not ( n8663 , n7809 );
not ( n8664 , n24 );
not ( n8665 , n8298 );
or ( n8666 , n8664 , n8665 );
nand ( n8667 , n8666 , n7377 );
not ( n8668 , n8667 );
or ( n8669 , n8663 , n8668 );
not ( n8670 , n24 );
and ( n8671 , n8670 , n7376 );
nor ( n8672 , n8671 , n8627 );
nand ( n8673 , n8669 , n8672 );
nand ( n8674 , n8673 , n3082 , n8631 );
and ( n8675 , n96 , n8627 );
and ( n8676 , n724 , n8625 );
nor ( n8677 , n8675 , n8676 );
nand ( n8678 , n24 , n8390 );
and ( n8679 , n8678 , n7377 );
nor ( n8680 , n8679 , n295 );
nand ( n8681 , n7806 , n8680 );
nand ( n8682 , n24 , n8356 );
and ( n8683 , n7377 , n8682 );
nor ( n8684 , n8683 , n1316 );
nand ( n8685 , n8644 , n8684 );
nand ( n8686 , n8677 , n8681 , n7596 , n8685 );
nand ( n8687 , n42 , n6761 , n8686 );
and ( n8688 , n8662 , n8674 , n8687 );
and ( n8689 , n8641 , n8653 , n8688 );
nor ( n8690 , n1371 , n2791 );
not ( n8691 , n8644 );
not ( n8692 , n24 );
or ( n8693 , n8692 , n7538 );
nand ( n8694 , n8693 , n7377 );
not ( n8695 , n8694 );
or ( n8696 , n8691 , n8695 );
nand ( n8697 , n8696 , n8626 );
and ( n8698 , n8690 , n8697 );
not ( n8699 , n24 );
or ( n8700 , n8699 , n8547 );
nand ( n8701 , n8700 , n7377 );
and ( n8702 , n8644 , n8701 );
nor ( n8703 , n8702 , n8625 );
or ( n8704 , n8703 , n1371 , n2450 );
not ( n8705 , n8644 );
not ( n8706 , n24 );
not ( n8707 , n8510 );
or ( n8708 , n8706 , n8707 );
nand ( n8709 , n8708 , n7377 );
not ( n8710 , n8709 );
or ( n8711 , n8705 , n8710 );
nand ( n8712 , n8711 , n8626 );
nand ( n8713 , n570 , n8712 );
or ( n8714 , n2303 , n18 , n8713 );
nand ( n8715 , n8704 , n8714 );
not ( n8716 , n42 );
nand ( n8717 , n1406 , n435 );
not ( n8718 , n24 );
not ( n8719 , n7728 );
or ( n8720 , n8718 , n8719 );
nand ( n8721 , n8720 , n7377 );
and ( n8722 , n8644 , n8721 );
nor ( n8723 , n8722 , n8625 );
nor ( n8724 , n8716 , n8717 , n8723 , n14 );
nor ( n8725 , n8698 , n8715 , n8724 );
not ( n8726 , n8644 );
not ( n8727 , n96 );
not ( n8728 , n24 );
not ( n8729 , n8469 );
or ( n8730 , n8728 , n8729 );
nand ( n8731 , n8730 , n7377 );
not ( n8732 , n8731 );
or ( n8733 , n8727 , n8732 );
not ( n8734 , n24 );
not ( n8735 , n8478 );
or ( n8736 , n8734 , n8735 );
nand ( n8737 , n8736 , n7377 );
and ( n8738 , n724 , n8737 );
nor ( n8739 , n8738 , n7957 );
nand ( n8740 , n8733 , n8739 );
not ( n8741 , n8740 );
or ( n8742 , n8726 , n8741 );
not ( n8743 , n3435 );
nor ( n8744 , n8743 , n8626 );
nor ( n8745 , n8744 , n7957 );
nand ( n8746 , n8742 , n8745 );
and ( n8747 , n42 , n2746 , n8746 );
not ( n8748 , n24 );
not ( n8749 , n8748 );
not ( n8750 , n8535 );
and ( n8751 , n8749 , n8750 );
nor ( n8752 , n8751 , n7376 );
or ( n8753 , n8645 , n8752 );
nand ( n8754 , n8753 , n8626 );
and ( n8755 , n42 , n1924 , n8754 );
nor ( n8756 , n8747 , n8755 );
and ( n8757 , n7806 , n7647 );
nor ( n8758 , n8757 , n8627 );
not ( n8759 , n8758 );
and ( n8760 , n3413 , n8759 );
and ( n8761 , n8644 , n7437 );
nor ( n8762 , n8761 , n8625 );
or ( n8763 , n3305 , n8762 );
not ( n8764 , n7704 );
nand ( n8765 , n8763 , n8764 );
nor ( n8766 , n8760 , n8765 );
not ( n8767 , n8644 );
not ( n8768 , n24 );
not ( n8769 , n7939 );
or ( n8770 , n8768 , n8769 );
nand ( n8771 , n8770 , n7377 );
not ( n8772 , n8771 );
or ( n8773 , n8767 , n8772 );
nand ( n8774 , n8773 , n8626 );
and ( n8775 , n2489 , n8774 );
and ( n8776 , n8644 , n7546 );
nor ( n8777 , n8776 , n8625 );
not ( n8778 , n8777 );
and ( n8779 , n3281 , n8778 );
nor ( n8780 , n8775 , n8779 );
and ( n8781 , n3345 , n7415 );
not ( n8782 , n7787 );
nor ( n8783 , n8781 , n8782 );
and ( n8784 , n8766 , n8780 , n8783 , n7788 );
nand ( n8785 , n2385 , n2818 );
and ( n8786 , n8644 , n7682 );
nor ( n8787 , n8786 , n8625 );
or ( n8788 , n8785 , n8787 );
and ( n8789 , n8644 , n7514 );
nor ( n8790 , n8789 , n8625 );
or ( n8791 , n7516 , n8790 );
nand ( n8792 , n8788 , n8791 );
nor ( n8793 , n8792 , n7417 , n7563 );
and ( n8794 , n8644 , n7692 );
nor ( n8795 , n8794 , n8625 );
not ( n8796 , n8795 );
and ( n8797 , n2418 , n8796 );
and ( n8798 , n8644 , n7378 );
nor ( n8799 , n8798 , n8625 );
not ( n8800 , n8799 );
and ( n8801 , n2463 , n8800 );
nor ( n8802 , n8797 , n8801 );
not ( n8803 , n2436 );
nor ( n8804 , n2303 , n8803 );
not ( n8805 , n8804 );
or ( n8806 , n8645 , n7782 );
nor ( n8807 , n8744 , n7557 );
nand ( n8808 , n3352 , n8625 );
nand ( n8809 , n8806 , n8807 , n8808 );
not ( n8810 , n8809 );
or ( n8811 , n8805 , n8810 );
not ( n8812 , n19 );
not ( n8813 , n8644 );
not ( n8814 , n7624 );
or ( n8815 , n8813 , n8814 );
nand ( n8816 , n8815 , n8745 );
nand ( n8817 , n8812 , n2461 , n8816 );
nand ( n8818 , n8811 , n8817 );
nor ( n8819 , n7652 , n8818 );
nand ( n8820 , n8784 , n8793 , n8802 , n8819 );
and ( n8821 , n18 , n8820 );
not ( n8822 , n24 );
not ( n8823 , n8413 );
or ( n8824 , n8822 , n8823 );
nand ( n8825 , n8824 , n7377 );
not ( n8826 , n8825 );
or ( n8827 , n8826 , n8645 );
nand ( n8828 , n8827 , n8626 );
and ( n8829 , n42 , n1787 , n8828 );
nor ( n8830 , n8821 , n8829 );
nand ( n8831 , n8689 , n8725 , n8756 , n8830 );
not ( n8832 , n8831 );
or ( n8833 , n8607 , n8832 );
nand ( n8834 , n8771 , n7380 , n2489 );
nand ( n8835 , n8833 , n8834 );
not ( n8836 , n8835 );
not ( n8837 , n3797 );
not ( n8838 , n8837 );
not ( n8839 , n8831 );
or ( n8840 , n8838 , n8839 );
not ( n8841 , n3800 );
nor ( n8842 , n18 , n8841 );
not ( n8843 , n7788 );
and ( n8844 , n3221 , n8721 );
and ( n8845 , n2418 , n8701 );
nor ( n8846 , n8844 , n8845 );
nand ( n8847 , n8846 , n7698 , n8783 );
not ( n8848 , n3281 );
not ( n8849 , n8694 );
or ( n8850 , n8848 , n8849 );
nand ( n8851 , n8850 , n7703 );
nor ( n8852 , n8843 , n8847 , n8851 , n7562 );
and ( n8853 , n2489 , n8658 );
or ( n8854 , n7516 , n8647 );
not ( n8855 , n8613 );
or ( n8856 , n2551 , n8855 );
nand ( n8857 , n8854 , n8856 );
nor ( n8858 , n8853 , n8857 , n7417 );
and ( n8859 , n2463 , n8709 );
nor ( n8860 , n8859 , n7559 , n7652 );
not ( n8861 , n8530 );
not ( n8862 , n8752 );
and ( n8863 , n8861 , n8862 );
not ( n8864 , n8804 );
not ( n8865 , n8680 );
not ( n8866 , n8684 );
nand ( n8867 , n8865 , n7596 , n8866 );
not ( n8868 , n8867 );
or ( n8869 , n8864 , n8868 );
nand ( n8870 , n453 , n8740 );
or ( n8871 , n2303 , n8870 );
not ( n8872 , n8785 );
and ( n8873 , n8872 , n8667 );
and ( n8874 , n3413 , n8825 );
nor ( n8875 , n8873 , n8874 );
nand ( n8876 , n8869 , n8871 , n8875 );
nor ( n8877 , n8863 , n8876 );
nand ( n8878 , n8852 , n8858 , n8860 , n8877 );
nand ( n8879 , n8842 , n3521 , n8878 );
nand ( n8880 , n8840 , n8879 );
not ( n8881 , n8880 );
nand ( n8882 , n7650 , n8606 , n8836 , n8881 );
nand ( n8883 , n7296 , n2506 , n8882 );
not ( n8884 , n4249 );
and ( n8885 , n2299 , n3569 , n4183 );
not ( n8886 , n8885 );
nor ( n8887 , n8884 , n8886 );
and ( n8888 , n914 , n8658 );
or ( n8889 , n912 , n7817 );
nor ( n8890 , n3454 , n7558 );
not ( n8891 , n8890 );
nand ( n8892 , n8889 , n8891 );
nor ( n8893 , n8888 , n8892 );
or ( n8894 , n963 , n8752 );
and ( n8895 , n909 , n8667 );
not ( n8896 , n8567 );
and ( n8897 , n8896 , n8721 );
nor ( n8898 , n8895 , n8897 );
and ( n8899 , n2440 , n8867 );
nor ( n8900 , n2387 , n434 );
and ( n8901 , n8900 , n8613 );
nor ( n8902 , n8899 , n8901 );
nand ( n8903 , n8893 , n8894 , n8898 , n8902 );
and ( n8904 , n3121 , n8903 );
nor ( n8905 , n3236 , n2190 );
and ( n8906 , n590 , n8905 );
and ( n8907 , n8906 , n7647 );
nor ( n8908 , n8904 , n8907 );
or ( n8909 , n20 , n7951 , n8227 );
not ( n8910 , n8012 );
nand ( n8911 , n8909 , n8910 );
and ( n8912 , n520 , n7682 );
and ( n8913 , n590 , n8771 );
nor ( n8914 , n8912 , n8913 );
or ( n8915 , n3288 , n8914 );
nor ( n8916 , n7949 , n438 );
nand ( n8917 , n1547 , n8916 );
or ( n8918 , n8917 , n8149 );
or ( n8919 , n7953 , n7817 );
nand ( n8920 , n8915 , n8918 , n8919 );
or ( n8921 , n8241 , n632 , n7953 );
not ( n8922 , n8602 );
not ( n8923 , n8900 );
or ( n8924 , n8528 , n8922 , n8923 );
nand ( n8925 , n8921 , n8924 );
and ( n8926 , n8602 , n8890 );
nor ( n8927 , n3311 , n7558 );
and ( n8928 , n13 , n8927 );
nor ( n8929 , n8926 , n8928 );
nor ( n8930 , n7949 , n8251 );
and ( n8931 , n8191 , n2193 , n8930 );
nor ( n8932 , n3346 , n7558 );
not ( n8933 , n8932 );
nand ( n8934 , n3256 , n7557 );
nand ( n8935 , n8933 , n8934 );
and ( n8936 , n7950 , n8935 );
nor ( n8937 , n8931 , n8936 );
and ( n8938 , n7514 , n520 , n8905 );
nor ( n8939 , n3236 , n438 );
and ( n8940 , n7692 , n1561 , n8939 );
nor ( n8941 , n8938 , n8940 );
and ( n8942 , n8197 , n1561 , n8916 );
nor ( n8943 , n8273 , n7953 , n521 );
nor ( n8944 , n8942 , n8943 );
nand ( n8945 , n8929 , n8937 , n8941 , n8944 );
nor ( n8946 , n8911 , n8920 , n8925 , n8945 );
and ( n8947 , n8541 , n8602 , n942 );
not ( n8948 , n8185 );
or ( n8949 , n8948 , n7949 , n2196 );
not ( n8950 , n438 );
nand ( n8951 , n8602 , n8950 , n2382 , n8561 );
nand ( n8952 , n8949 , n8951 );
nor ( n8953 , n8947 , n8952 );
nor ( n8954 , n13 , n1989 );
and ( n8955 , n8954 , n7437 );
nand ( n8956 , n7378 , n3250 , n570 );
and ( n8957 , n3250 , n8935 );
not ( n8958 , n13 );
and ( n8959 , n8958 , n8927 );
nor ( n8960 , n8957 , n8959 );
nand ( n8961 , n8956 , n8960 );
or ( n8962 , n3238 , n7783 );
and ( n8963 , n7546 , n1547 , n8939 );
not ( n8964 , n3292 );
not ( n8965 , n8905 );
and ( n8966 , n8964 , n8965 );
nor ( n8967 , n8966 , n7817 );
nor ( n8968 , n8963 , n8967 );
not ( n8969 , n20 );
nand ( n8970 , n8969 , n3237 , n7624 );
nand ( n8971 , n8962 , n8968 , n8970 );
nor ( n8972 , n8955 , n8961 , n8971 );
and ( n8973 , n8908 , n8946 , n8953 , n8972 );
and ( n8974 , n766 , n8825 );
and ( n8975 , n8125 , n8701 );
not ( n8976 , n3264 );
and ( n8977 , n8976 , n8694 );
nor ( n8978 , n8974 , n8975 , n8977 );
not ( n8979 , n8647 );
and ( n8980 , n584 , n8979 );
not ( n8981 , n19 );
and ( n8982 , n8981 , n1407 );
nor ( n8983 , n8982 , n20 , n7558 );
nor ( n8984 , n8980 , n8983 );
nand ( n8985 , n570 , n8709 );
nand ( n8986 , n8978 , n8984 , n8985 , n8870 );
and ( n8987 , n3121 , n8986 );
not ( n8988 , n8930 );
nor ( n8989 , n8266 , n912 , n8988 );
nor ( n8990 , n8987 , n8989 );
nand ( n8991 , n8338 , n908 , n8602 );
or ( n8992 , n6283 , n8550 );
not ( n8993 , n8514 );
and ( n8994 , n570 , n8993 );
nor ( n8995 , n8994 , n8932 );
not ( n8996 , n8976 );
not ( n8997 , n8584 );
or ( n8998 , n8996 , n8997 );
nand ( n8999 , n8998 , n8934 );
not ( n9000 , n2195 );
not ( n9001 , n8441 );
or ( n9002 , n9000 , n9001 );
not ( n9003 , n8494 );
or ( n9004 , n841 , n9003 );
nand ( n9005 , n9002 , n9004 );
nor ( n9006 , n8999 , n9005 );
nand ( n9007 , n8992 , n8995 , n9006 );
or ( n9008 , n8393 , n9007 );
nand ( n9009 , n9008 , n8602 );
nand ( n9010 , n8973 , n8990 , n8991 , n9009 );
nand ( n9011 , n8887 , n7794 , n9010 );
and ( n9012 , n4250 , n4223 );
nand ( n9013 , n2508 , n9012 , n8831 );
not ( n9014 , n6 );
nor ( n9015 , n2506 , n7 );
and ( n9016 , n9015 , n7793 );
nand ( n9017 , n9014 , n8885 , n18 , n9016 );
not ( n9018 , n9017 );
nand ( n9019 , n9018 , n8950 );
or ( n9020 , n9019 , n1548 , n8777 );
or ( n9021 , n8799 , n571 , n9017 );
nand ( n9022 , n9020 , n9021 );
or ( n9023 , n8795 , n6283 , n9017 );
not ( n9024 , n1592 );
nand ( n9025 , n8885 , n4249 , n7793 );
or ( n9026 , n8762 , n9024 , n9025 );
nand ( n9027 , n9023 , n9026 );
nor ( n9028 , n9022 , n9027 );
not ( n9029 , n9025 );
not ( n9030 , n8927 );
not ( n9031 , n9030 );
and ( n9032 , n9029 , n9031 );
not ( n9033 , n8935 );
nor ( n9034 , n9033 , n9017 );
nor ( n9035 , n9032 , n9034 );
not ( n9036 , n9035 );
nand ( n9037 , n18 , n19 );
nor ( n9038 , n20 , n9037 );
not ( n9039 , n9038 );
nor ( n9040 , n7817 , n9039 , n9025 );
nor ( n9041 , n9036 , n9040 );
nand ( n9042 , n24 , n4261 );
not ( n9043 , n18 );
nand ( n9044 , n9043 , n9015 , n7793 );
nor ( n9045 , n9044 , n6 , n8886 );
and ( n9046 , n8900 , n8629 );
nor ( n9047 , n9046 , n8892 , n8661 );
not ( n9048 , n8723 );
nand ( n9049 , n9048 , n8896 );
not ( n9050 , n2441 );
and ( n9051 , n9050 , n8686 );
and ( n9052 , n909 , n8673 );
and ( n9053 , n942 , n8754 );
nor ( n9054 , n9051 , n9052 , n9053 );
nand ( n9055 , n9047 , n9049 , n9054 );
and ( n9056 , n9045 , n9055 );
nand ( n9057 , n3242 , n7793 );
nand ( n9058 , n4249 , n8885 , n520 );
or ( n9059 , n8787 , n9057 , n9058 );
not ( n9060 , n7817 );
nand ( n9061 , n4249 , n9060 );
or ( n9062 , n9061 , n8886 , n9057 );
nand ( n9063 , n9059 , n9062 );
nand ( n9064 , n9038 , n7793 );
nor ( n9065 , n8790 , n9064 , n9058 );
nor ( n9066 , n9056 , n9063 , n9065 );
nand ( n9067 , n9028 , n9041 , n9042 , n9066 );
and ( n9068 , n3425 , n8809 );
and ( n9069 , n2009 , n8816 );
nor ( n9070 , n9068 , n9069 );
or ( n9071 , n9025 , n9070 );
or ( n9072 , n6283 , n8703 );
and ( n9073 , n766 , n8828 );
not ( n9074 , n8713 );
nor ( n9075 , n9073 , n8983 , n9074 );
and ( n9076 , n453 , n8746 );
and ( n9077 , n8976 , n8697 );
and ( n9078 , n584 , n8649 );
nor ( n9079 , n9076 , n9077 , n9078 );
nand ( n9080 , n9072 , n9075 , n9079 );
and ( n9081 , n9045 , n9080 );
nand ( n9082 , n590 , n4249 , n8885 );
nor ( n9083 , n8758 , n9064 , n9082 );
nor ( n9084 , n9081 , n9083 );
not ( n9085 , n9057 );
not ( n9086 , n9082 );
nand ( n9087 , n9085 , n8774 , n9086 );
not ( n9088 , n4323 );
not ( n9089 , n9088 );
nand ( n9090 , n24 , n9089 , n7389 );
nand ( n9091 , n9090 , n7368 , n7812 );
and ( n9092 , n8900 , n9091 );
and ( n9093 , n2392 , n7555 );
nor ( n9094 , n9092 , n9093 );
or ( n9095 , n3928 , n9094 );
nand ( n9096 , n3090 , n3787 );
nand ( n9097 , n450 , n9091 );
and ( n9098 , n7414 , n9097 );
or ( n9099 , n9096 , n9098 );
not ( n9100 , n9096 );
not ( n9101 , n9091 );
or ( n9102 , n2228 , n9101 );
nand ( n9103 , n9102 , n7556 );
not ( n9104 , n9103 );
not ( n9105 , n9104 );
and ( n9106 , n9100 , n9105 );
not ( n9107 , n3747 );
nand ( n9108 , n3242 , n9107 );
and ( n9109 , n3435 , n9091 );
nor ( n9110 , n9109 , n7957 );
nor ( n9111 , n9108 , n9110 );
nor ( n9112 , n9106 , n9111 );
nand ( n9113 , n9095 , n9099 , n9112 );
not ( n9114 , n7396 );
not ( n9115 , n3748 );
or ( n9116 , n9114 , n3516 , n9115 );
not ( n9117 , n3748 );
or ( n9118 , n9117 , n7558 );
nand ( n9119 , n9116 , n9118 );
not ( n9120 , n646 );
nor ( n9121 , n16 , n9120 );
not ( n9122 , n9121 );
or ( n9123 , n9098 , n9122 , n3928 );
not ( n9124 , n8265 );
or ( n9125 , n3748 , n9024 , n9124 );
nand ( n9126 , n9123 , n9125 );
nor ( n9127 , n9113 , n9119 , n9126 );
or ( n9128 , n3089 , n9104 );
or ( n9129 , n912 , n9110 );
or ( n9130 , n2067 , n9098 );
nand ( n9131 , n9128 , n9129 , n9130 );
nand ( n9132 , n450 , n7821 );
nor ( n9133 , n8016 , n9122 , n9132 );
or ( n9134 , n8923 , n8527 );
or ( n9135 , n3090 , n9121 );
not ( n9136 , n9098 );
nand ( n9137 , n9135 , n9136 );
nand ( n9138 , n9134 , n9137 );
nor ( n9139 , n9131 , n9133 , n9138 );
and ( n9140 , n2066 , n9103 );
or ( n9141 , n963 , n8540 );
nand ( n9142 , n9141 , n9094 );
nor ( n9143 , n9140 , n9142 );
nor ( n9144 , n2067 , n7822 );
and ( n9145 , n8377 , n450 , n9144 );
not ( n9146 , n9132 );
and ( n9147 , n8335 , n3090 , n9146 );
nor ( n9148 , n9145 , n9147 );
and ( n9149 , n8368 , n2229 , n9144 );
nand ( n9150 , n2229 , n7821 );
not ( n9151 , n9150 );
and ( n9152 , n8325 , n3090 , n9151 );
nor ( n9153 , n9149 , n9152 );
nand ( n9154 , n9139 , n9143 , n9148 , n9153 );
and ( n9155 , n3990 , n9154 );
or ( n9156 , n8275 , n9096 , n9150 );
nand ( n9157 , n2066 , n3787 );
or ( n9158 , n8243 , n9157 , n9150 );
nand ( n9159 , n9156 , n9158 );
not ( n9160 , n8240 );
nor ( n9161 , n8923 , n3928 , n9160 );
nor ( n9162 , n9155 , n9159 , n9161 );
nor ( n9163 , n7651 , n9150 );
not ( n9164 , n9163 );
or ( n9165 , n9164 , n8204 );
nor ( n9166 , n2186 , n7822 );
nand ( n9167 , n2229 , n9166 );
or ( n9168 , n9167 , n8231 );
nor ( n9169 , n571 , n7822 );
not ( n9170 , n9169 );
or ( n9171 , n9170 , n8156 );
nand ( n9172 , n9165 , n9168 , n9171 );
not ( n9173 , n9172 );
nand ( n9174 , n454 , n9136 );
not ( n9175 , n9174 );
nor ( n9176 , n1931 , n9098 );
nor ( n9177 , n7651 , n9104 );
nor ( n9178 , n9176 , n9177 );
nand ( n9179 , n3146 , n7555 );
nand ( n9180 , n8976 , n9091 );
nand ( n9181 , n9178 , n9179 , n9180 );
nor ( n9182 , n1931 , n9132 );
not ( n9183 , n9182 );
or ( n9184 , n9183 , n8123 );
nand ( n9185 , n2458 , n9136 );
nand ( n9186 , n9184 , n9185 );
nor ( n9187 , n2186 , n9104 );
nor ( n9188 , n9175 , n9181 , n9186 , n9187 );
and ( n9189 , n8976 , n8148 );
nor ( n9190 , n3176 , n9110 );
not ( n9191 , n9190 );
nor ( n9192 , n7651 , n9132 );
nand ( n9193 , n9192 , n8116 );
nand ( n9194 , n9191 , n9193 );
nand ( n9195 , n450 , n9166 );
nor ( n9196 , n9195 , n8095 );
nor ( n9197 , n9189 , n9194 , n9196 );
nand ( n9198 , n9173 , n9188 , n9197 );
and ( n9199 , n3787 , n9198 );
nand ( n9200 , n9121 , n3787 , n9146 , n8020 );
not ( n9201 , n9096 );
nand ( n9202 , n9201 , n7913 , n9146 );
nand ( n9203 , n9200 , n9202 );
nor ( n9204 , n9199 , n9203 );
not ( n9205 , n8583 );
and ( n9206 , n8976 , n9205 );
and ( n9207 , n9182 , n8522 );
nor ( n9208 , n9206 , n9207 );
nand ( n9209 , n9185 , n9208 , n9179 , n9180 );
nor ( n9210 , n9209 , n9176 , n9177 );
or ( n9211 , n9195 , n8496 );
nand ( n9212 , n9211 , n9174 );
nor ( n9213 , n9212 , n9187 , n9190 );
and ( n9214 , n9192 , n8427 );
and ( n9215 , n9169 , n8506 );
nor ( n9216 , n9214 , n9215 );
not ( n9217 , n9167 );
not ( n9218 , n8587 );
and ( n9219 , n9217 , n9218 );
and ( n9220 , n9163 , n8436 );
nor ( n9221 , n9219 , n9220 );
nand ( n9222 , n9210 , n9213 , n9216 , n9221 );
and ( n9223 , n3990 , n9222 );
and ( n9224 , n9098 , n9104 );
nor ( n9225 , n9224 , n9157 );
nor ( n9226 , n8259 , n9157 , n9132 );
nor ( n9227 , n9223 , n9225 , n9226 );
nand ( n9228 , n9127 , n9162 , n9204 , n9227 );
nand ( n9229 , n4258 , n9228 );
nand ( n9230 , n9071 , n9084 , n9087 , n9229 );
nor ( n9231 , n9067 , n9230 );
nand ( n9232 , n8883 , n9011 , n9013 , n9231 );
nand ( n9233 , n25 , n34 );
not ( n9234 , n30 );
nor ( n9235 , n27 , n166 );
nand ( n9236 , n9234 , n9235 );
not ( n9237 , n9236 );
not ( n9238 , n9237 );
nand ( n9239 , n25 , n9238 );
not ( n9240 , n26 );
not ( n9241 , n9240 );
not ( n9242 , n4385 );
not ( n9243 , n30 );
nand ( n9244 , n9243 , n7300 );
nand ( n9245 , n9242 , n9244 );
not ( n9246 , n9245 );
not ( n9247 , n9246 );
or ( n9248 , n9241 , n9247 );
nand ( n9249 , n9248 , n234 );
and ( n9250 , n9239 , n9249 );
nand ( n9251 , n9233 , n9250 );
not ( n9252 , n9251 );
or ( n9253 , n17 , n9252 );
not ( n9254 , n22 );
or ( n9255 , n9254 , n9233 );
and ( n9256 , n22 , n25 );
not ( n9257 , n9256 );
not ( n9258 , n28 );
not ( n9259 , n391 );
or ( n9260 , n9258 , n9259 );
nand ( n9261 , n9260 , n7301 );
not ( n9262 , n9261 );
or ( n9263 , n9257 , n9262 );
not ( n9264 , n25 );
nand ( n9265 , n9264 , n22 );
not ( n9266 , n26 );
not ( n9267 , n28 );
nand ( n9268 , n9267 , n9244 );
not ( n9269 , n9268 );
nand ( n9270 , n9266 , n9269 );
not ( n9271 , n9270 );
or ( n9272 , n9265 , n9271 );
nand ( n9273 , n9263 , n9272 );
not ( n9274 , n9273 );
nand ( n9275 , n9255 , n9274 );
not ( n9276 , n9275 );
or ( n9277 , n692 , n9276 );
and ( n9278 , n31 , n274 );
and ( n9279 , n21 , n9278 );
nor ( n9280 , n9279 , n15 );
and ( n9281 , n17 , n9280 );
not ( n9282 , n17 );
nand ( n9283 , n21 , n31 , n15 , n7374 );
and ( n9284 , n9282 , n9283 );
nor ( n9285 , n9281 , n9284 );
nand ( n9286 , n9253 , n9277 , n9285 );
and ( n9287 , n16 , n9038 , n9286 );
nand ( n9288 , n2191 , n3437 );
and ( n9289 , n9024 , n9288 );
and ( n9290 , n42 , n4323 );
nor ( n9291 , n9289 , n21 , n9290 );
nor ( n9292 , n9287 , n9291 );
not ( n9293 , n25 );
and ( n9294 , n7332 , n4493 );
buf ( n9295 , n9294 );
not ( n9296 , n9295 );
not ( n9297 , n9296 );
or ( n9298 , n9293 , n9297 );
not ( n9299 , n26 );
not ( n9300 , n4288 );
not ( n9301 , n9300 );
nand ( n9302 , n9301 , n9244 );
not ( n9303 , n9302 );
and ( n9304 , n9299 , n9303 );
nor ( n9305 , n9304 , n25 );
not ( n9306 , n9305 );
nand ( n9307 , n9298 , n9306 );
not ( n9308 , n9307 );
or ( n9309 , n21 , n9308 );
and ( n9310 , n21 , n462 , n9307 );
not ( n9311 , n21 );
nor ( n9312 , n9311 , n23 );
nand ( n9313 , n31 , n9312 );
or ( n9314 , n9313 , n9274 );
nor ( n9315 , n22 , n9313 );
not ( n9316 , n9315 );
or ( n9317 , n9316 , n9250 );
not ( n9318 , n21 );
not ( n9319 , n22 );
nand ( n9320 , n9319 , n23 );
or ( n9321 , n9318 , n9320 );
not ( n9322 , n9321 );
not ( n9323 , n9296 );
not ( n9324 , n9323 );
and ( n9325 , n9322 , n9324 );
not ( n9326 , n21 );
or ( n9327 , n9326 , n100 );
not ( n9328 , n4290 );
not ( n9329 , n9328 );
nor ( n9330 , n9327 , n9329 );
nor ( n9331 , n9325 , n9330 );
nand ( n9332 , n9314 , n9317 , n9331 );
nor ( n9333 , n9310 , n9332 );
nand ( n9334 , n9309 , n9333 );
and ( n9335 , n1592 , n9334 );
or ( n9336 , n17 , n9250 );
or ( n9337 , n692 , n9274 );
nand ( n9338 , n9336 , n9337 , n9285 );
and ( n9339 , n1975 , n9338 );
nor ( n9340 , n9335 , n9339 );
nor ( n9341 , n2244 , n7651 );
not ( n9342 , n35 );
and ( n9343 , n22 , n9342 );
nor ( n9344 , n25 , n32 );
nand ( n9345 , n26 , n9344 );
buf ( n9346 , n9344 );
and ( n9347 , n232 , n9268 );
nand ( n9348 , n9346 , n9347 );
nand ( n9349 , n9345 , n9348 );
nand ( n9350 , n9343 , n9349 );
nand ( n9351 , n22 , n549 );
nand ( n9352 , n234 , n9270 );
or ( n9353 , n9351 , n9352 );
not ( n9354 , n9343 );
nor ( n9355 , n32 , n220 );
not ( n9356 , n9355 );
or ( n9357 , n9354 , n9356 );
nand ( n9358 , n9256 , n549 );
nand ( n9359 , n9357 , n9358 );
not ( n9360 , n33 );
not ( n9361 , n9360 );
not ( n9362 , n655 );
or ( n9363 , n9361 , n9362 );
not ( n9364 , n34 );
nand ( n9365 , n33 , n9261 );
nand ( n9366 , n9364 , n9365 );
not ( n9367 , n9366 );
nand ( n9368 , n9363 , n9367 );
nand ( n9369 , n9359 , n9368 );
and ( n9370 , n9350 , n9353 , n9369 );
or ( n9371 , n15 , n9370 );
not ( n9372 , n9280 );
nand ( n9373 , n9371 , n9372 );
and ( n9374 , n9341 , n18 , n9373 );
nor ( n9375 , n22 , n35 );
not ( n9376 , n9375 );
or ( n9377 , n7491 , n9376 );
not ( n9378 , n25 );
nor ( n9379 , n9378 , n22 );
not ( n9380 , n9379 );
nand ( n9381 , n9377 , n9380 );
not ( n9382 , n33 );
not ( n9383 , n9382 );
not ( n9384 , n7448 );
not ( n9385 , n9384 );
or ( n9386 , n9383 , n9385 );
nor ( n9387 , n34 , n9238 );
nand ( n9388 , n9386 , n9387 );
nand ( n9389 , n9381 , n9388 );
nand ( n9390 , n232 , n9245 );
not ( n9391 , n9390 );
not ( n9392 , n9346 );
nor ( n9393 , n9392 , n9376 );
nand ( n9394 , n9391 , n9393 );
not ( n9395 , n22 );
and ( n9396 , n9395 , n549 );
nand ( n9397 , n234 , n9245 );
nor ( n9398 , n26 , n9397 );
and ( n9399 , n9396 , n9398 );
nor ( n9400 , n22 , n25 );
nand ( n9401 , n26 , n9400 );
not ( n9402 , n9401 );
nor ( n9403 , n9399 , n9402 );
and ( n9404 , n9389 , n9394 , n9403 );
or ( n9405 , n17 , n9404 );
not ( n9406 , n9284 );
nand ( n9407 , n9405 , n9406 );
not ( n9408 , n14 );
not ( n9409 , n18 );
nor ( n9410 , n9408 , n9409 );
and ( n9411 , n9407 , n9410 , n2458 );
nor ( n9412 , n9374 , n9411 );
not ( n9413 , n9288 );
not ( n9414 , n21 );
not ( n9415 , n9414 );
not ( n9416 , n25 );
nand ( n9417 , n4512 , n9294 );
buf ( n9418 , n9417 );
not ( n9419 , n9418 );
or ( n9420 , n9416 , n9419 );
nand ( n9421 , n9420 , n9306 );
not ( n9422 , n9421 );
not ( n9423 , n9422 );
not ( n9424 , n9423 );
or ( n9425 , n9415 , n9424 );
not ( n9426 , n23 );
nand ( n9427 , n9426 , n5063 );
not ( n9428 , n9427 );
and ( n9429 , n9428 , n9421 );
and ( n9430 , n9315 , n9251 );
nor ( n9431 , n9429 , n9430 );
not ( n9432 , n9313 );
and ( n9433 , n9432 , n9275 );
not ( n9434 , n9418 );
or ( n9435 , n9321 , n9434 );
not ( n9436 , n9330 );
nand ( n9437 , n9435 , n9436 );
nor ( n9438 , n9433 , n9437 );
and ( n9439 , n9431 , n9438 );
nand ( n9440 , n9425 , n9439 );
and ( n9441 , n9413 , n9440 );
nor ( n9442 , n16 , n1581 );
not ( n9443 , n21 );
nand ( n9444 , n9443 , n2229 );
nor ( n9445 , n9444 , n9290 );
and ( n9446 , n9442 , n9445 );
nor ( n9447 , n9441 , n9446 );
and ( n9448 , n9292 , n9340 , n9412 , n9447 );
and ( n9449 , n25 , n549 );
not ( n9450 , n33 );
not ( n9451 , n9450 );
not ( n9452 , n34 );
nand ( n9453 , n9452 , n4618 , n9294 );
not ( n9454 , n9453 );
or ( n9455 , n9451 , n9454 );
nand ( n9456 , n33 , n9417 );
nand ( n9457 , n9455 , n9456 );
nand ( n9458 , n9449 , n9457 );
not ( n9459 , n9305 );
or ( n9460 , n550 , n9459 );
not ( n9461 , n35 );
not ( n9462 , n9355 );
not ( n9463 , n9457 );
or ( n9464 , n9462 , n9463 );
nand ( n9465 , n234 , n4372 , n9302 );
nand ( n9466 , n9345 , n9465 );
not ( n9467 , n9466 );
nand ( n9468 , n9464 , n9467 );
nand ( n9469 , n9461 , n9468 );
nand ( n9470 , n9458 , n9460 , n9469 );
not ( n9471 , n9470 );
or ( n9472 , n9427 , n9471 );
or ( n9473 , n9313 , n9370 );
not ( n9474 , n35 );
not ( n9475 , n9327 );
nand ( n9476 , n9474 , n9475 );
not ( n9477 , n32 );
nand ( n9478 , n9477 , n4607 );
nand ( n9479 , n32 , n9328 );
nand ( n9480 , n9478 , n4346 , n9479 );
not ( n9481 , n9480 );
or ( n9482 , n9476 , n9481 );
nand ( n9483 , n21 , n23 );
nand ( n9484 , n22 , n35 );
nor ( n9485 , n9483 , n9484 );
not ( n9486 , n9329 );
nand ( n9487 , n9485 , n9486 );
nand ( n9488 , n9482 , n9487 );
or ( n9489 , n9313 , n9404 );
nand ( n9490 , n9322 , n9457 );
nand ( n9491 , n9489 , n9490 );
nor ( n9492 , n9488 , n9491 );
nand ( n9493 , n9472 , n9473 , n9492 );
and ( n9494 , n9493 , n2385 , n2866 );
not ( n9495 , n18 );
nor ( n9496 , n9495 , n2303 );
not ( n9497 , n31 );
nand ( n9498 , n9497 , n15 );
not ( n9499 , n9498 );
and ( n9500 , n9499 , n8619 );
not ( n9501 , n9500 );
nand ( n9502 , n37 , n9245 );
not ( n9503 , n9502 );
nand ( n9504 , n9503 , n9393 );
not ( n9505 , n9380 );
not ( n9506 , n37 );
not ( n9507 , n32 );
nand ( n9508 , n9506 , n9507 , n9375 );
not ( n9509 , n9508 );
or ( n9510 , n9505 , n9509 );
not ( n9511 , n9236 );
not ( n9512 , n9511 );
not ( n9513 , n33 );
nand ( n9514 , n9512 , n9513 );
nand ( n9515 , n34 , n9514 );
nand ( n9516 , n33 , n9238 );
not ( n9517 , n33 );
nand ( n9518 , n36 , n9237 );
nand ( n9519 , n9517 , n9518 );
nand ( n9520 , n9515 , n9516 , n9519 );
nand ( n9521 , n9510 , n9520 );
nand ( n9522 , n9504 , n9403 , n9521 );
not ( n9523 , n9522 );
or ( n9524 , n17 , n9523 );
nand ( n9525 , n9524 , n9406 );
nor ( n9526 , n9501 , n9525 );
nor ( n9527 , n9417 , n4460 );
or ( n9528 , n33 , n9527 );
nand ( n9529 , n9528 , n9456 );
nand ( n9530 , n9449 , n9529 );
not ( n9531 , n35 );
nor ( n9532 , n32 , n477 );
not ( n9533 , n9532 );
not ( n9534 , n9529 );
or ( n9535 , n9533 , n9534 );
nand ( n9536 , n234 , n606 , n9302 );
nand ( n9537 , n9345 , n9536 );
not ( n9538 , n9537 );
nand ( n9539 , n9535 , n9538 );
nand ( n9540 , n9531 , n9539 );
nand ( n9541 , n9530 , n9460 , n9540 );
buf ( n9542 , n9541 );
not ( n9543 , n9542 );
not ( n9544 , n9543 );
not ( n9545 , n9544 );
not ( n9546 , n9428 );
not ( n9547 , n9542 );
or ( n9548 , n9546 , n9547 );
not ( n9549 , n9476 );
or ( n9550 , n32 , n4441 );
nand ( n9551 , n9479 , n9550 , n4438 );
nand ( n9552 , n9549 , n9551 );
and ( n9553 , n9487 , n9552 );
nand ( n9554 , n9548 , n9553 );
nand ( n9555 , n9322 , n9529 );
and ( n9556 , n9343 , n9532 );
not ( n9557 , n9358 );
nor ( n9558 , n9556 , n9557 );
not ( n9559 , n33 );
not ( n9560 , n397 );
not ( n9561 , n9560 );
and ( n9562 , n9559 , n9561 );
nor ( n9563 , n9562 , n9366 );
or ( n9564 , n9558 , n9563 );
nor ( n9565 , n232 , n9269 );
nand ( n9566 , n9346 , n9565 );
nand ( n9567 , n9345 , n9566 );
nand ( n9568 , n9343 , n9567 );
nand ( n9569 , n9564 , n9568 , n9353 );
or ( n9570 , n9522 , n9569 );
nand ( n9571 , n9570 , n9432 );
nand ( n9572 , n9555 , n9571 );
nor ( n9573 , n9554 , n9572 );
and ( n9574 , n9526 , n9545 , n9573 );
or ( n9575 , n2065 , n9573 );
not ( n9576 , n14 );
and ( n9577 , n9576 , n9525 );
or ( n9578 , n15 , n2344 );
not ( n9579 , n9578 );
and ( n9580 , n9579 , n9569 );
nor ( n9581 , n9577 , n9580 );
not ( n9582 , n21 );
nand ( n9583 , n9582 , n2345 );
or ( n9584 , n9278 , n9578 );
and ( n9585 , n9583 , n9584 );
nand ( n9586 , n9575 , n9581 , n9585 );
nand ( n9587 , n2458 , n9586 );
nor ( n9588 , n9574 , n9587 );
and ( n9589 , n9496 , n9588 );
nor ( n9590 , n9494 , n9589 );
nor ( n9591 , n1984 , n2384 );
not ( n9592 , n33 );
not ( n9593 , n9592 );
nand ( n9594 , n7333 , n4559 , n4363 );
not ( n9595 , n9594 );
or ( n9596 , n9593 , n9595 );
nand ( n9597 , n33 , n9296 );
nand ( n9598 , n9596 , n9597 );
nand ( n9599 , n9449 , n9598 );
not ( n9600 , n35 );
not ( n9601 , n9355 );
not ( n9602 , n9598 );
or ( n9603 , n9601 , n9602 );
nand ( n9604 , n9603 , n9467 );
nand ( n9605 , n9600 , n9604 );
nand ( n9606 , n9599 , n9460 , n9605 );
not ( n9607 , n9606 );
or ( n9608 , n9427 , n9607 );
nand ( n9609 , n9322 , n9598 );
nand ( n9610 , n9608 , n9609 );
not ( n9611 , n9249 );
not ( n9612 , n9611 );
not ( n9613 , n9612 );
nand ( n9614 , n7448 , n9237 );
not ( n9615 , n9614 );
or ( n9616 , n33 , n9615 );
nand ( n9617 , n9616 , n9516 );
nand ( n9618 , n25 , n9617 );
not ( n9619 , n9618 );
or ( n9620 , n9613 , n9619 );
nand ( n9621 , n9620 , n9396 );
not ( n9622 , n32 );
not ( n9623 , n9622 );
not ( n9624 , n9618 );
not ( n9625 , n9624 );
or ( n9626 , n9623 , n9625 );
and ( n9627 , n7492 , n9617 );
not ( n9628 , n26 );
not ( n9629 , n9628 );
not ( n9630 , n9390 );
or ( n9631 , n9629 , n9630 );
nand ( n9632 , n9631 , n9346 );
not ( n9633 , n9632 );
nor ( n9634 , n9627 , n9633 );
nand ( n9635 , n9626 , n9634 );
nand ( n9636 , n9375 , n9635 );
and ( n9637 , n9621 , n9636 );
nand ( n9638 , n160 , n9261 );
not ( n9639 , n9638 );
not ( n9640 , n34 );
not ( n9641 , n9261 );
or ( n9642 , n9640 , n9641 );
buf ( n9643 , n175 );
nand ( n9644 , n9642 , n9643 );
not ( n9645 , n9644 );
nand ( n9646 , n7450 , n9645 );
nand ( n9647 , n203 , n9646 );
not ( n9648 , n9647 );
or ( n9649 , n9639 , n9648 );
not ( n9650 , n32 );
nand ( n9651 , n9649 , n9650 );
or ( n9652 , n26 , n9347 );
not ( n9653 , n9346 );
not ( n9654 , n9653 );
nand ( n9655 , n9652 , n9654 );
not ( n9656 , n9365 );
not ( n9657 , n33 );
nand ( n9658 , n9657 , n9646 );
not ( n9659 , n9658 );
or ( n9660 , n9656 , n9659 );
not ( n9661 , n7492 );
not ( n9662 , n9661 );
nand ( n9663 , n9660 , n9662 );
nand ( n9664 , n9651 , n9655 , n9663 );
and ( n9665 , n9343 , n9664 );
and ( n9666 , n9352 , n9638 );
and ( n9667 , n9666 , n9647 );
nor ( n9668 , n9667 , n9351 );
nor ( n9669 , n9665 , n9668 );
and ( n9670 , n9637 , n9669 );
nor ( n9671 , n9670 , n9313 );
nor ( n9672 , n9610 , n9488 , n9671 );
not ( n9673 , n9672 );
and ( n9674 , n2229 , n9673 );
or ( n9675 , n17 , n9637 );
nand ( n9676 , n9675 , n9406 );
and ( n9677 , n14 , n9676 );
nor ( n9678 , n9674 , n9677 , n9445 );
or ( n9679 , n15 , n9669 );
not ( n9680 , n9372 );
not ( n9681 , n9680 );
not ( n9682 , n9681 );
not ( n9683 , n9682 );
nand ( n9684 , n9679 , n9683 );
and ( n9685 , n2245 , n9684 );
not ( n9686 , n9444 );
and ( n9687 , n9686 , n9606 );
nor ( n9688 , n9685 , n9687 );
not ( n9689 , n33 );
not ( n9690 , n34 );
not ( n9691 , n9690 );
not ( n9692 , n4457 );
or ( n9693 , n9691 , n9692 );
nand ( n9694 , n9693 , n9294 );
nand ( n9695 , n9689 , n9694 );
nand ( n9696 , n9597 , n9695 );
nand ( n9697 , n9449 , n9696 );
not ( n9698 , n35 );
not ( n9699 , n9532 );
not ( n9700 , n9696 );
or ( n9701 , n9699 , n9700 );
not ( n9702 , n9537 );
nand ( n9703 , n9701 , n9702 );
nand ( n9704 , n9698 , n9703 );
nand ( n9705 , n9460 , n9697 , n9704 );
not ( n9706 , n9705 );
not ( n9707 , n9706 );
not ( n9708 , n9707 );
nand ( n9709 , n9322 , n9696 );
and ( n9710 , n9709 , n9553 );
nand ( n9711 , n9428 , n9707 );
not ( n9712 , n7533 );
not ( n9713 , n9712 );
not ( n9714 , n9713 );
not ( n9715 , n33 );
not ( n9716 , n9715 );
not ( n9717 , n384 );
nand ( n9718 , n9717 , n9511 );
not ( n9719 , n9718 );
or ( n9720 , n9716 , n9719 );
nand ( n9721 , n9720 , n9516 );
and ( n9722 , n9714 , n9721 );
not ( n9723 , n32 );
not ( n9724 , n9723 );
not ( n9725 , n9718 );
or ( n9726 , n200 , n9725 );
not ( n9727 , n9237 );
nand ( n9728 , n158 , n9727 );
nand ( n9729 , n9726 , n9728 );
not ( n9730 , n9729 );
or ( n9731 , n9724 , n9730 );
not ( n9732 , n26 );
not ( n9733 , n9732 );
not ( n9734 , n9502 );
or ( n9735 , n9733 , n9734 );
nand ( n9736 , n9735 , n9346 );
nand ( n9737 , n9731 , n9736 );
nor ( n9738 , n9722 , n9737 );
or ( n9739 , n9376 , n9738 );
or ( n9740 , n9611 , n9729 );
nand ( n9741 , n9740 , n9396 );
nand ( n9742 , n9739 , n9741 );
not ( n9743 , n9742 );
not ( n9744 , n9743 );
not ( n9745 , n9343 );
not ( n9746 , n9638 );
not ( n9747 , n385 );
not ( n9748 , n9747 );
nand ( n9749 , n9748 , n9645 );
nand ( n9750 , n203 , n9749 );
not ( n9751 , n9750 );
or ( n9752 , n9746 , n9751 );
not ( n9753 , n32 );
nand ( n9754 , n9752 , n9753 );
or ( n9755 , n26 , n9565 );
nand ( n9756 , n9755 , n9654 );
not ( n9757 , n9365 );
not ( n9758 , n33 );
nand ( n9759 , n9758 , n9749 );
not ( n9760 , n9759 );
or ( n9761 , n9757 , n9760 );
not ( n9762 , n9713 );
nand ( n9763 , n9761 , n9762 );
nand ( n9764 , n9754 , n9756 , n9763 );
not ( n9765 , n9764 );
or ( n9766 , n9745 , n9765 );
not ( n9767 , n9666 );
not ( n9768 , n9750 );
or ( n9769 , n9767 , n9768 );
not ( n9770 , n9351 );
nand ( n9771 , n9769 , n9770 );
nand ( n9772 , n9766 , n9771 );
or ( n9773 , n9744 , n9772 );
nand ( n9774 , n9773 , n9432 );
nand ( n9775 , n9710 , n9711 , n9774 );
not ( n9776 , n9775 );
and ( n9777 , n9708 , n9776 );
and ( n9778 , n9579 , n9772 );
not ( n9779 , n14 );
not ( n9780 , n9779 );
or ( n9781 , n17 , n9743 );
nand ( n9782 , n9781 , n9406 );
not ( n9783 , n9782 );
or ( n9784 , n9780 , n9783 );
nand ( n9785 , n9784 , n9585 );
nor ( n9786 , n9778 , n9785 );
nor ( n9787 , n9777 , n9786 );
not ( n9788 , n9787 );
nand ( n9789 , n450 , n9775 );
or ( n9790 , n9501 , n9782 );
nand ( n9791 , n9786 , n9789 );
nand ( n9792 , n9790 , n9791 );
nand ( n9793 , n9788 , n9789 , n9792 );
and ( n9794 , n42 , n9793 );
buf ( n9795 , n9791 );
and ( n9796 , n2303 , n9795 );
nor ( n9797 , n9794 , n9796 );
nand ( n9798 , n9678 , n9688 , n9797 );
and ( n9799 , n9591 , n9798 );
not ( n9800 , n18 );
nor ( n9801 , n9800 , n9587 );
and ( n9802 , n2303 , n9801 );
nor ( n9803 , n9799 , n9802 );
and ( n9804 , n9590 , n9803 );
not ( n9805 , n16 );
nand ( n9806 , n9805 , n2879 );
not ( n9807 , n17 );
or ( n9808 , n32 , n476 );
not ( n9809 , n22 );
nand ( n9810 , n9808 , n9809 );
nor ( n9811 , n9810 , n9725 );
not ( n9812 , n9400 );
nor ( n9813 , n32 , n9812 );
not ( n9814 , n9813 );
not ( n9815 , n9503 );
or ( n9816 , n9814 , n9815 );
nand ( n9817 , n9816 , n9401 );
nor ( n9818 , n9811 , n9817 );
and ( n9819 , n25 , n7533 );
nor ( n9820 , n9819 , n1383 );
or ( n9821 , n9818 , n9820 );
not ( n9822 , n22 );
not ( n9823 , n9397 );
nand ( n9824 , n9822 , n1382 , n9823 );
nand ( n9825 , n9821 , n9824 );
and ( n9826 , n9807 , n9825 );
nor ( n9827 , n9826 , n9284 );
or ( n9828 , n14 , n9827 );
nand ( n9829 , n22 , n1382 );
not ( n9830 , n32 );
nand ( n9831 , n9830 , n379 );
and ( n9832 , n25 , n9831 );
nor ( n9833 , n9829 , n9832 );
and ( n9834 , n22 , n232 );
and ( n9835 , n22 , n32 );
nor ( n9836 , n9834 , n9835 );
not ( n9837 , n9836 );
not ( n9838 , n9749 );
not ( n9839 , n9838 );
and ( n9840 , n9837 , n9839 );
nor ( n9841 , n32 , n9265 );
and ( n9842 , n9841 , n9565 );
nor ( n9843 , n9840 , n9842 );
nand ( n9844 , n22 , n9832 );
not ( n9845 , n9844 );
not ( n9846 , n9838 );
and ( n9847 , n9845 , n9846 );
nand ( n9848 , n22 , n26 );
nor ( n9849 , n9848 , n9832 );
nor ( n9850 , n9847 , n9849 );
and ( n9851 , n9843 , n9850 );
or ( n9852 , n9833 , n9851 );
not ( n9853 , n7491 );
or ( n9854 , n26 , n9853 );
nand ( n9855 , n9854 , n25 );
nor ( n9856 , n25 , n9269 );
nand ( n9857 , n9855 , n9835 , n9856 );
nand ( n9858 , n9852 , n9857 );
nand ( n9859 , n9579 , n9858 );
nand ( n9860 , n9828 , n9585 , n9859 );
and ( n9861 , n9501 , n9860 );
not ( n9862 , n350 );
not ( n9863 , n9694 );
and ( n9864 , n7383 , n9863 );
not ( n9865 , n32 );
nor ( n9866 , n9864 , n9865 );
not ( n9867 , n9866 );
or ( n9868 , n9862 , n9867 );
not ( n9869 , n26 );
nand ( n9870 , n32 , n9869 , n234 , n9302 );
not ( n9871 , n9870 );
not ( n9872 , n9532 );
not ( n9873 , n9694 );
or ( n9874 , n9872 , n9873 );
not ( n9875 , n9537 );
nand ( n9876 , n9874 , n9875 );
nor ( n9877 , n9871 , n9876 );
nand ( n9878 , n9868 , n9877 );
not ( n9879 , n9878 );
and ( n9880 , n9827 , n9879 );
nand ( n9881 , n9322 , n9694 );
and ( n9882 , n9428 , n9878 );
and ( n9883 , n9432 , n9825 );
nor ( n9884 , n9882 , n9883 );
and ( n9885 , n9881 , n9884 );
nand ( n9886 , n9475 , n9551 );
nand ( n9887 , n9432 , n9858 );
nand ( n9888 , n9885 , n9886 , n9887 );
and ( n9889 , n450 , n9888 );
nor ( n9890 , n9889 , n9860 );
nor ( n9891 , n9880 , n9890 );
not ( n9892 , n9860 );
and ( n9893 , n2065 , n9892 );
not ( n9894 , n9888 );
nor ( n9895 , n9893 , n9894 );
nor ( n9896 , n9861 , n9891 , n9895 );
or ( n9897 , n9806 , n9896 );
nand ( n9898 , n2816 , n2229 );
not ( n9899 , n33 );
not ( n9900 , n9295 );
nand ( n9901 , n9899 , n9900 );
nand ( n9902 , n33 , n9594 );
and ( n9903 , n9901 , n9902 );
not ( n9904 , n9903 );
and ( n9905 , n25 , n256 );
nand ( n9906 , n9904 , n9905 );
or ( n9907 , n255 , n9306 );
not ( n9908 , n9355 );
or ( n9909 , n9908 , n9903 );
nand ( n9910 , n9909 , n9467 );
nand ( n9911 , n35 , n9910 );
nand ( n9912 , n9906 , n9907 , n9911 );
and ( n9913 , n9428 , n9912 );
nor ( n9914 , n9321 , n9903 );
nor ( n9915 , n9913 , n9914 );
and ( n9916 , n9485 , n9480 );
not ( n9917 , n9486 );
nor ( n9918 , n9476 , n9917 );
nor ( n9919 , n9916 , n9918 );
not ( n9920 , n22 );
and ( n9921 , n35 , n9920 );
and ( n9922 , n33 , n9614 );
not ( n9923 , n9514 );
nor ( n9924 , n9922 , n9923 );
nor ( n9925 , n234 , n9924 );
not ( n9926 , n9925 );
or ( n9927 , n32 , n9926 );
or ( n9928 , n9661 , n9924 );
nand ( n9929 , n9927 , n9928 , n9632 );
and ( n9930 , n9921 , n9929 );
or ( n9931 , n9925 , n9611 );
nor ( n9932 , n22 , n255 );
nand ( n9933 , n9931 , n9932 );
not ( n9934 , n9933 );
nor ( n9935 , n9930 , n9934 );
not ( n9936 , n9935 );
not ( n9937 , n161 );
nand ( n9938 , n9937 , n9646 );
not ( n9939 , n9261 );
not ( n9940 , n9939 );
not ( n9941 , n33 );
nand ( n9942 , n9940 , n9941 );
not ( n9943 , n9942 );
nand ( n9944 , n25 , n9943 );
and ( n9945 , n9938 , n9352 , n9944 );
not ( n9946 , n22 );
nor ( n9947 , n9946 , n255 );
not ( n9948 , n9947 );
nor ( n9949 , n9945 , n9948 );
not ( n9950 , n202 );
nand ( n9951 , n9950 , n9261 );
not ( n9952 , n9951 );
not ( n9953 , n9938 );
or ( n9954 , n9952 , n9953 );
not ( n9955 , n32 );
nand ( n9956 , n9954 , n9955 );
not ( n9957 , n9942 );
nand ( n9958 , n33 , n9646 );
not ( n9959 , n9958 );
or ( n9960 , n9957 , n9959 );
nand ( n9961 , n9960 , n9662 );
and ( n9962 , n9956 , n9655 , n9961 );
nor ( n9963 , n9962 , n9484 );
nor ( n9964 , n9949 , n9963 );
not ( n9965 , n9964 );
or ( n9966 , n9936 , n9965 );
nand ( n9967 , n9966 , n9432 );
nand ( n9968 , n9915 , n9919 , n9967 );
not ( n9969 , n9968 );
or ( n9970 , n9898 , n9969 );
not ( n9971 , n16 );
not ( n9972 , n19 );
nand ( n9973 , n9972 , n9686 );
nor ( n9974 , n9971 , n9973 );
not ( n9975 , n9912 );
not ( n9976 , n9975 );
and ( n9977 , n9974 , n9976 );
not ( n9978 , n2126 );
nor ( n9979 , n9327 , n9481 );
and ( n9980 , n9978 , n9979 );
not ( n9981 , n14 );
or ( n9982 , n17 , n9981 , n1407 );
nand ( n9983 , n9432 , n830 );
nand ( n9984 , n9982 , n9983 );
nand ( n9985 , n4351 , n1382 );
not ( n9986 , n9985 );
not ( n9987 , n32 );
and ( n9988 , n9987 , n7577 );
nor ( n9989 , n9988 , n22 );
and ( n9990 , n9989 , n9614 );
and ( n9991 , n9813 , n9391 );
nor ( n9992 , n9991 , n9402 );
not ( n9993 , n9992 );
nor ( n9994 , n9990 , n9993 );
or ( n9995 , n9986 , n9994 );
nand ( n9996 , n9995 , n9824 );
and ( n9997 , n9984 , n9996 );
not ( n9998 , n6679 );
nand ( n9999 , n92 , n9998 );
and ( n10000 , n9999 , n9983 );
not ( n10001 , n9835 );
nand ( n10002 , n22 , n7576 );
not ( n10003 , n9646 );
or ( n10004 , n10002 , n10003 );
and ( n10005 , n9841 , n9347 );
nor ( n10006 , n10005 , n9849 );
nand ( n10007 , n10004 , n10006 );
and ( n10008 , n10001 , n10007 );
not ( n10009 , n10001 );
not ( n10010 , n10002 );
or ( n10011 , n10009 , n10010 );
nand ( n10012 , n10011 , n9646 );
and ( n10013 , n10006 , n10012 );
or ( n10014 , n4606 , n10013 );
nand ( n10015 , n10014 , n9857 );
nor ( n10016 , n10008 , n10015 );
nor ( n10017 , n10000 , n10016 );
nor ( n10018 , n9980 , n9997 , n10017 );
not ( n10019 , n9594 );
not ( n10020 , n10019 );
nand ( n10021 , n10020 , n9322 , n2127 );
and ( n10022 , n3299 , n9284 );
and ( n10023 , n9998 , n9680 );
nor ( n10024 , n10022 , n10023 );
nand ( n10025 , n10018 , n10021 , n10024 );
nor ( n10026 , n9977 , n10025 );
nand ( n10027 , n9970 , n10026 );
nand ( n10028 , n16 , n2879 );
not ( n10029 , n33 );
or ( n10030 , n10029 , n9863 );
nand ( n10031 , n10030 , n9901 );
nand ( n10032 , n9322 , n10031 );
and ( n10033 , n9485 , n9551 );
nor ( n10034 , n10033 , n9918 );
and ( n10035 , n10032 , n10034 );
nand ( n10036 , n9905 , n10031 );
not ( n10037 , n9532 );
not ( n10038 , n10031 );
or ( n10039 , n10037 , n10038 );
nand ( n10040 , n10039 , n9538 );
nand ( n10041 , n35 , n10040 );
nand ( n10042 , n10036 , n9907 , n10041 );
nand ( n10043 , n9428 , n10042 );
not ( n10044 , n9932 );
or ( n10045 , n234 , n9514 );
nand ( n10046 , n158 , n9718 );
nand ( n10047 , n10045 , n9249 , n10046 );
not ( n10048 , n10047 );
or ( n10049 , n10044 , n10048 );
not ( n10050 , n9921 );
nand ( n10051 , n199 , n9238 );
not ( n10052 , n10051 );
not ( n10053 , n10046 );
or ( n10054 , n10052 , n10053 );
not ( n10055 , n32 );
nand ( n10056 , n10054 , n10055 );
not ( n10057 , n33 );
not ( n10058 , n9718 );
or ( n10059 , n10057 , n10058 );
nand ( n10060 , n10059 , n9514 );
nand ( n10061 , n9712 , n10060 );
nand ( n10062 , n10056 , n9736 , n10061 );
not ( n10063 , n10062 );
or ( n10064 , n10050 , n10063 );
nand ( n10065 , n10049 , n10064 );
not ( n10066 , n10065 );
not ( n10067 , n10066 );
not ( n10068 , n9947 );
not ( n10069 , n161 );
nand ( n10070 , n10069 , n9749 );
nand ( n10071 , n10070 , n9352 , n9944 );
not ( n10072 , n10071 );
or ( n10073 , n10068 , n10072 );
not ( n10074 , n9484 );
not ( n10075 , n9951 );
not ( n10076 , n10070 );
or ( n10077 , n10075 , n10076 );
not ( n10078 , n32 );
nand ( n10079 , n10077 , n10078 );
not ( n10080 , n9942 );
nand ( n10081 , n33 , n9749 );
not ( n10082 , n10081 );
or ( n10083 , n10080 , n10082 );
nand ( n10084 , n10083 , n9762 );
nand ( n10085 , n10079 , n9756 , n10084 );
nand ( n10086 , n10074 , n10085 );
nand ( n10087 , n10073 , n10086 );
not ( n10088 , n10087 );
not ( n10089 , n10088 );
or ( n10090 , n10067 , n10089 );
nand ( n10091 , n10090 , n9432 );
nand ( n10092 , n10035 , n10043 , n10091 );
or ( n10093 , n9501 , n10092 );
not ( n10094 , n14 );
or ( n10095 , n17 , n10066 );
nand ( n10096 , n10095 , n9406 );
and ( n10097 , n10094 , n10096 );
or ( n10098 , n9578 , n10088 );
nand ( n10099 , n10098 , n9585 );
nor ( n10100 , n10097 , n10099 );
not ( n10101 , n10100 );
nand ( n10102 , n10093 , n10101 );
nand ( n10103 , n450 , n10092 );
or ( n10104 , n10042 , n10096 );
nand ( n10105 , n10100 , n10103 );
nand ( n10106 , n10104 , n10105 );
and ( n10107 , n10102 , n10103 , n10106 );
or ( n10108 , n10028 , n10107 );
and ( n10109 , n2816 , n10105 );
not ( n10110 , n9890 );
and ( n10111 , n2332 , n10110 );
nor ( n10112 , n10109 , n10111 );
or ( n10113 , n42 , n10112 );
nand ( n10114 , n2816 , n9445 );
not ( n10115 , n10114 );
not ( n10116 , n9290 );
nor ( n10117 , n21 , n1995 );
and ( n10118 , n14 , n10116 , n10117 );
nor ( n10119 , n10115 , n10118 );
nand ( n10120 , n10108 , n10113 , n10119 );
nor ( n10121 , n10027 , n10120 );
not ( n10122 , n1937 );
nand ( n10123 , n9428 , n10122 );
not ( n10124 , n7369 );
not ( n10125 , n10124 );
not ( n10126 , n10019 );
or ( n10127 , n10125 , n10126 );
nand ( n10128 , n10127 , n32 );
not ( n10129 , n10128 );
nand ( n10130 , n7521 , n10129 );
and ( n10131 , n9355 , n9594 );
nor ( n10132 , n10131 , n9466 );
and ( n10133 , n10130 , n9870 , n10132 );
nor ( n10134 , n10123 , n10133 );
or ( n10135 , n17 , n9935 );
nand ( n10136 , n10135 , n9406 );
nand ( n10137 , n6835 , n10136 );
not ( n10138 , n10137 );
not ( n10139 , n9978 );
nor ( n10140 , n21 , n10139 );
not ( n10141 , n10140 );
not ( n10142 , n10133 );
not ( n10143 , n10142 );
or ( n10144 , n10141 , n10143 );
not ( n10145 , n16 );
not ( n10146 , n6678 );
nor ( n10147 , n10145 , n10146 );
or ( n10148 , n15 , n9964 );
nand ( n10149 , n10148 , n9683 );
nand ( n10150 , n10147 , n10149 );
nand ( n10151 , n10144 , n10150 );
nor ( n10152 , n10134 , n10138 , n10151 );
nand ( n10153 , n9897 , n10121 , n10152 );
and ( n10154 , n1582 , n10153 );
buf ( n10155 , n2534 );
not ( n10156 , n9313 );
nor ( n10157 , n10001 , n4351 );
not ( n10158 , n7302 );
and ( n10159 , n171 , n10158 );
nand ( n10160 , n9747 , n10159 );
and ( n10161 , n10157 , n10160 );
not ( n10162 , n9829 );
nand ( n10163 , n10162 , n9856 );
not ( n10164 , n10163 );
and ( n10165 , n26 , n10160 );
nor ( n10166 , n10165 , n7524 );
nand ( n10167 , n9355 , n10160 );
and ( n10168 , n10166 , n9348 , n10167 );
not ( n10169 , n22 );
nor ( n10170 , n10168 , n10169 );
nor ( n10171 , n10161 , n10164 , n10170 );
not ( n10172 , n10171 );
and ( n10173 , n10156 , n10172 );
nor ( n10174 , n10173 , n9979 );
not ( n10175 , n4618 );
not ( n10176 , n10175 );
not ( n10177 , n34 );
nand ( n10178 , n10176 , n10177 , n9295 );
not ( n10179 , n10178 );
not ( n10180 , n10179 );
nand ( n10181 , n9322 , n10180 );
and ( n10182 , n9355 , n10178 );
not ( n10183 , n9302 );
nor ( n10184 , n10183 , n32 , n37 , n25 );
nor ( n10185 , n10182 , n10184 );
nand ( n10186 , n25 , n10179 );
nand ( n10187 , n4334 , n10186 );
and ( n10188 , n10185 , n9870 , n10187 );
nand ( n10189 , n26 , n10186 );
not ( n10190 , n4351 );
not ( n10191 , n26 );
nand ( n10192 , n10191 , n10180 );
not ( n10193 , n10192 );
not ( n10194 , n10189 );
or ( n10195 , n10193 , n10194 );
nand ( n10196 , n10195 , n32 );
and ( n10197 , n10187 , n10185 );
nand ( n10198 , n10196 , n10197 );
nand ( n10199 , n10190 , n10198 );
nand ( n10200 , n10188 , n10189 , n10199 );
and ( n10201 , n9428 , n10200 );
not ( n10202 , n9985 );
not ( n10203 , n9387 );
or ( n10204 , n7451 , n10203 );
nand ( n10205 , n10204 , n9989 );
nand ( n10206 , n9992 , n10205 );
not ( n10207 , n10206 );
or ( n10208 , n10202 , n10207 );
nand ( n10209 , n10208 , n9824 );
and ( n10210 , n9432 , n10209 );
nor ( n10211 , n10201 , n10210 );
nand ( n10212 , n10174 , n10181 , n10211 );
and ( n10213 , n10155 , n10212 );
not ( n10214 , n17 );
and ( n10215 , n9384 , n9237 );
nor ( n10216 , n10215 , n9810 );
nor ( n10217 , n10216 , n9817 );
or ( n10218 , n9820 , n10217 );
nand ( n10219 , n10218 , n9824 );
and ( n10220 , n10214 , n10219 );
nor ( n10221 , n10220 , n9284 );
or ( n10222 , n14 , n10221 );
nand ( n10223 , n7449 , n10159 );
nand ( n10224 , n10157 , n10223 );
not ( n10225 , n26 );
not ( n10226 , n10223 );
or ( n10227 , n10225 , n10226 );
nand ( n10228 , n10227 , n7383 );
not ( n10229 , n10228 );
nand ( n10230 , n9532 , n10223 );
nand ( n10231 , n10229 , n9566 , n10230 );
nand ( n10232 , n22 , n10231 );
and ( n10233 , n10224 , n10163 , n10232 );
or ( n10234 , n10233 , n9578 );
nand ( n10235 , n10222 , n10234 , n9585 );
nand ( n10236 , n9501 , n10235 );
or ( n10237 , n450 , n10235 );
or ( n10238 , n9313 , n10233 );
not ( n10239 , n9886 );
buf ( n10240 , n7334 );
not ( n10241 , n10240 );
nand ( n10242 , n10241 , n4678 );
not ( n10243 , n10242 );
nor ( n10244 , n9321 , n10243 );
nor ( n10245 , n10239 , n10244 );
not ( n10246 , n7521 );
buf ( n10247 , n10124 );
and ( n10248 , n10247 , n10243 );
not ( n10249 , n32 );
nor ( n10250 , n10248 , n10249 );
not ( n10251 , n10250 );
or ( n10252 , n10246 , n10251 );
not ( n10253 , n9532 );
not ( n10254 , n10242 );
or ( n10255 , n10253 , n10254 );
nand ( n10256 , n10255 , n9702 );
nor ( n10257 , n9871 , n10256 );
nand ( n10258 , n10252 , n10257 );
and ( n10259 , n9428 , n10258 );
and ( n10260 , n9432 , n10219 );
nor ( n10261 , n10259 , n10260 );
nand ( n10262 , n10238 , n10245 , n10261 );
nand ( n10263 , n10237 , n10262 );
not ( n10264 , n10221 );
not ( n10265 , n10258 );
not ( n10266 , n10265 );
or ( n10267 , n10264 , n10266 );
not ( n10268 , n450 );
not ( n10269 , n10262 );
or ( n10270 , n10268 , n10269 );
not ( n10271 , n10235 );
nand ( n10272 , n10270 , n10271 );
nand ( n10273 , n10267 , n10272 );
and ( n10274 , n10236 , n10263 , n10273 );
or ( n10275 , n9806 , n10274 );
not ( n10276 , n7491 );
and ( n10277 , n9921 , n10276 );
nor ( n10278 , n10277 , n9379 );
not ( n10279 , n33 );
nor ( n10280 , n10279 , n34 );
and ( n10281 , n36 , n10280 );
nor ( n10282 , n10281 , n10203 );
or ( n10283 , n10278 , n10282 );
nor ( n10284 , n10050 , n9653 );
nand ( n10285 , n9391 , n10284 );
and ( n10286 , n9932 , n9398 );
nor ( n10287 , n10286 , n9402 );
and ( n10288 , n10283 , n10285 , n10287 );
nand ( n10289 , n10074 , n9349 );
not ( n10290 , n9352 );
nand ( n10291 , n9947 , n10290 );
not ( n10292 , n9256 );
nor ( n10293 , n10292 , n255 );
nor ( n10294 , n9484 , n9908 );
or ( n10295 , n10293 , n10294 );
not ( n10296 , n33 );
not ( n10297 , n655 );
or ( n10298 , n10296 , n10297 );
not ( n10299 , n34 );
nand ( n10300 , n10299 , n9942 );
not ( n10301 , n10300 );
nand ( n10302 , n10298 , n10301 );
nand ( n10303 , n10295 , n10302 );
and ( n10304 , n10289 , n10291 , n10303 );
and ( n10305 , n10288 , n10304 );
nor ( n10306 , n10305 , n9313 );
not ( n10307 , n33 );
not ( n10308 , n10178 );
or ( n10309 , n10307 , n10308 );
not ( n10310 , n33 );
nand ( n10311 , n10310 , n9418 );
nand ( n10312 , n10309 , n10311 );
nand ( n10313 , n9905 , n10312 );
not ( n10314 , n9355 );
not ( n10315 , n10312 );
or ( n10316 , n10314 , n10315 );
nand ( n10317 , n10316 , n9467 );
nand ( n10318 , n35 , n10317 );
nand ( n10319 , n10313 , n9907 , n10318 );
not ( n10320 , n10319 );
or ( n10321 , n9427 , n10320 );
nand ( n10322 , n9322 , n10312 );
nand ( n10323 , n10321 , n10322 , n9919 );
nor ( n10324 , n10306 , n10323 );
or ( n10325 , n9898 , n10324 );
not ( n10326 , n10028 );
not ( n10327 , n9428 );
not ( n10328 , n33 );
or ( n10329 , n10328 , n9527 );
nand ( n10330 , n10329 , n10311 );
nand ( n10331 , n9905 , n10330 );
not ( n10332 , n9532 );
not ( n10333 , n10330 );
or ( n10334 , n10332 , n10333 );
nand ( n10335 , n10334 , n9702 );
nand ( n10336 , n35 , n10335 );
nand ( n10337 , n10331 , n9907 , n10336 );
not ( n10338 , n10337 );
or ( n10339 , n10327 , n10338 );
nand ( n10340 , n10339 , n10034 );
nand ( n10341 , n9322 , n10330 );
and ( n10342 , n33 , n9518 );
not ( n10343 , n34 );
not ( n10344 , n9516 );
or ( n10345 , n10343 , n10344 );
nand ( n10346 , n10345 , n9514 );
nor ( n10347 , n10342 , n10346 );
not ( n10348 , n32 );
and ( n10349 , n232 , n10348 , n9921 );
nor ( n10350 , n10349 , n9379 );
or ( n10351 , n10347 , n10350 );
nand ( n10352 , n9503 , n10284 );
nand ( n10353 , n10351 , n10352 , n10287 );
and ( n10354 , n10074 , n9532 );
nor ( n10355 , n10354 , n10293 );
not ( n10356 , n33 );
nor ( n10357 , n10356 , n9560 );
nor ( n10358 , n10300 , n10357 );
or ( n10359 , n10355 , n10358 );
nand ( n10360 , n10074 , n9567 );
nand ( n10361 , n10359 , n10291 , n10360 );
or ( n10362 , n10353 , n10361 );
nand ( n10363 , n10362 , n9432 );
nand ( n10364 , n10341 , n10363 );
nor ( n10365 , n10340 , n10364 );
or ( n10366 , n2065 , n10365 );
not ( n10367 , n14 );
not ( n10368 , n17 );
and ( n10369 , n10368 , n10353 );
nor ( n10370 , n10369 , n9284 );
not ( n10371 , n10370 );
and ( n10372 , n10367 , n10371 );
and ( n10373 , n9579 , n10361 );
nor ( n10374 , n10372 , n10373 );
nand ( n10375 , n10366 , n10374 , n9585 );
not ( n10376 , n10337 );
nand ( n10377 , n9500 , n10370 , n10376 , n10365 );
nand ( n10378 , n10375 , n10377 );
not ( n10379 , n10378 );
and ( n10380 , n10326 , n10379 );
not ( n10381 , n16 );
nor ( n10382 , n19 , n42 );
not ( n10383 , n10382 );
nor ( n10384 , n10381 , n10383 );
and ( n10385 , n10384 , n10375 );
nor ( n10386 , n10380 , n10385 );
nand ( n10387 , n10275 , n10325 , n10386 );
not ( n10388 , n10140 );
not ( n10389 , n10200 );
or ( n10390 , n10388 , n10389 );
not ( n10391 , n16 );
nand ( n10392 , n10391 , n10382 );
not ( n10393 , n10272 );
or ( n10394 , n10392 , n10393 );
nand ( n10395 , n10390 , n10394 );
nor ( n10396 , n10213 , n10387 , n10395 );
or ( n10397 , n15 , n10304 );
nand ( n10398 , n10397 , n9372 );
and ( n10399 , n10147 , n10398 );
or ( n10400 , n17 , n10288 );
nand ( n10401 , n10400 , n9406 );
not ( n10402 , n10401 );
or ( n10403 , n6834 , n10402 );
nand ( n10404 , n10403 , n10119 );
nor ( n10405 , n10399 , n10404 );
not ( n10406 , n10320 );
not ( n10407 , n10406 );
not ( n10408 , n10407 );
and ( n10409 , n9974 , n10408 );
or ( n10410 , n15 , n10171 );
not ( n10411 , n9680 );
nand ( n10412 , n10410 , n10411 );
and ( n10413 , n9998 , n10412 );
not ( n10414 , n17 );
not ( n10415 , n10414 );
not ( n10416 , n10209 );
or ( n10417 , n10415 , n10416 );
nand ( n10418 , n10417 , n9406 );
and ( n10419 , n3299 , n10418 );
nor ( n10420 , n10409 , n10413 , n10419 );
nand ( n10421 , n10396 , n10405 , n10420 );
and ( n10422 , n309 , n10421 );
nor ( n10423 , n10154 , n10422 );
not ( n10424 , n18 );
not ( n10425 , n21 );
nand ( n10426 , n10425 , n570 , n10116 );
nor ( n10427 , n22 , n32 );
and ( n10428 , n10427 , n9251 );
not ( n10429 , n22 );
nand ( n10430 , n10429 , n32 );
not ( n10431 , n10430 );
not ( n10432 , n34 );
not ( n10433 , n7455 );
nand ( n10434 , n4885 , n10432 , n10124 , n10433 );
and ( n10435 , n10431 , n10434 );
nor ( n10436 , n10428 , n10435 );
or ( n10437 , n17 , n10436 );
and ( n10438 , n10001 , n9275 );
nand ( n10439 , n7383 , n9939 );
not ( n10440 , n10439 );
not ( n10441 , n34 );
nand ( n10442 , n10440 , n10441 );
and ( n10443 , n9835 , n10442 );
nor ( n10444 , n10438 , n10443 );
or ( n10445 , n692 , n10444 );
nand ( n10446 , n10437 , n10445 , n9285 );
and ( n10447 , n3345 , n10446 );
and ( n10448 , n2458 , n9445 );
nor ( n10449 , n10447 , n10448 );
not ( n10450 , n92 );
or ( n10451 , n9370 , n9835 );
not ( n10452 , n9368 );
or ( n10453 , n10001 , n10452 );
not ( n10454 , n9832 );
nand ( n10455 , n22 , n1104 , n10454 );
nand ( n10456 , n10451 , n10453 , n10455 );
not ( n10457 , n10456 );
or ( n10458 , n10450 , n10457 );
nand ( n10459 , n10458 , n9681 );
nand ( n10460 , n10459 , n2245 , n2458 );
not ( n10461 , n21 );
not ( n10462 , n10461 );
not ( n10463 , n32 );
nand ( n10464 , n10463 , n9421 );
not ( n10465 , n1387 );
nand ( n10466 , n32 , n9418 );
nand ( n10467 , n10464 , n10465 , n10466 );
not ( n10468 , n10467 );
or ( n10469 , n10462 , n10468 );
not ( n10470 , n32 );
or ( n10471 , n10470 , n2317 );
nand ( n10472 , n10471 , n10466 , n10464 );
and ( n10473 , n9428 , n10472 );
and ( n10474 , n10436 , n10444 );
nor ( n10475 , n10474 , n9313 );
not ( n10476 , n9437 );
not ( n10477 , n9483 );
nand ( n10478 , n10477 , n9835 );
nand ( n10479 , n10476 , n10478 );
nor ( n10480 , n10473 , n10475 , n10479 );
nand ( n10481 , n10469 , n10480 );
and ( n10482 , n782 , n10481 );
not ( n10483 , n17 );
not ( n10484 , n10483 );
or ( n10485 , n32 , n9404 );
or ( n10486 , n7371 , n9388 );
nand ( n10487 , n10486 , n10431 );
nand ( n10488 , n10485 , n10487 );
not ( n10489 , n10488 );
or ( n10490 , n10484 , n10489 );
nand ( n10491 , n10490 , n9406 );
and ( n10492 , n3251 , n10491 );
nor ( n10493 , n10482 , n10492 );
and ( n10494 , n10426 , n10449 , n10460 , n10493 );
nand ( n10495 , n32 , n9457 );
not ( n10496 , n32 );
nand ( n10497 , n10496 , n9470 );
nand ( n10498 , n10471 , n10495 , n9469 , n10497 );
nand ( n10499 , n2458 , n9686 , n10498 );
and ( n10500 , n10465 , n9540 );
nand ( n10501 , n32 , n9529 );
not ( n10502 , n32 );
nand ( n10503 , n10502 , n9541 );
nand ( n10504 , n10500 , n10501 , n10503 );
not ( n10505 , n10504 );
not ( n10506 , n10505 );
not ( n10507 , n450 );
not ( n10508 , n9343 );
not ( n10509 , n4721 );
not ( n10510 , n10509 );
or ( n10511 , n10508 , n10510 );
not ( n10512 , n35 );
or ( n10513 , n10512 , n9917 );
not ( n10514 , n32 );
nand ( n10515 , n10513 , n10514 );
nand ( n10516 , n22 , n10515 );
nand ( n10517 , n10511 , n10516 );
nand ( n10518 , n10477 , n10517 );
and ( n10519 , n10518 , n9555 );
and ( n10520 , n9428 , n10504 );
not ( n10521 , n32 );
and ( n10522 , n10521 , n9522 );
not ( n10523 , n9520 );
and ( n10524 , n10124 , n10523 );
nor ( n10525 , n10524 , n10430 );
nor ( n10526 , n10522 , n10525 );
and ( n10527 , n10001 , n9569 );
or ( n10528 , n10001 , n9563 );
nand ( n10529 , n10528 , n10455 );
nor ( n10530 , n10527 , n10529 );
and ( n10531 , n10526 , n10530 );
nor ( n10532 , n10531 , n9313 );
nor ( n10533 , n10520 , n10532 );
nand ( n10534 , n10519 , n10533 );
not ( n10535 , n10534 );
or ( n10536 , n10507 , n10535 );
not ( n10537 , n14 );
or ( n10538 , n17 , n10526 );
nand ( n10539 , n10538 , n9406 );
and ( n10540 , n10537 , n10539 );
or ( n10541 , n9578 , n10530 );
nand ( n10542 , n10541 , n9585 );
nor ( n10543 , n10540 , n10542 );
nand ( n10544 , n10536 , n10543 );
and ( n10545 , n10506 , n10544 );
nor ( n10546 , n9500 , n10543 );
nor ( n10547 , n10545 , n10546 );
and ( n10548 , n10539 , n10544 );
and ( n10549 , n10519 , n10533 );
and ( n10550 , n2065 , n10543 );
nor ( n10551 , n10549 , n10550 );
nor ( n10552 , n10548 , n10551 );
nand ( n10553 , n10547 , n10552 );
and ( n10554 , n10553 , n2385 , n2461 );
not ( n10555 , n9343 );
not ( n10556 , n4374 );
or ( n10557 , n10555 , n10556 );
nand ( n10558 , n10557 , n10516 );
nand ( n10559 , n10477 , n10558 );
and ( n10560 , n10559 , n9490 );
or ( n10561 , n10488 , n10456 );
nand ( n10562 , n10561 , n9432 );
and ( n10563 , n10465 , n10495 );
nand ( n10564 , n10563 , n9469 , n10497 );
nand ( n10565 , n9428 , n10564 );
nand ( n10566 , n10560 , n10562 , n10565 );
and ( n10567 , n10566 , n2229 , n2458 );
nor ( n10568 , n10554 , n10567 );
and ( n10569 , n10499 , n10568 );
nand ( n10570 , n10544 , n2385 , n2998 );
not ( n10571 , n20 );
not ( n10572 , n32 );
nor ( n10573 , n998 , n105 );
not ( n10574 , n10573 );
nor ( n10575 , n10572 , n10574 );
and ( n10576 , n10575 , n10228 );
not ( n10577 , n10223 );
nor ( n10578 , n10577 , n1383 , n10574 );
nor ( n10579 , n10576 , n10578 , n10244 );
or ( n10580 , n9313 , n10217 );
not ( n10581 , n32 );
and ( n10582 , n10581 , n9550 , n4438 );
nor ( n10583 , n10582 , n9327 );
not ( n10584 , n10583 );
nand ( n10585 , n10580 , n10584 );
not ( n10586 , n9428 );
not ( n10587 , n10250 );
not ( n10588 , n10256 );
nand ( n10589 , n10587 , n10588 );
not ( n10590 , n10589 );
or ( n10591 , n10586 , n10590 );
and ( n10592 , n234 , n9565 );
nor ( n10593 , n10592 , n10228 );
or ( n10594 , n32 , n10593 );
nand ( n10595 , n10594 , n10230 );
nand ( n10596 , n10573 , n10595 );
nand ( n10597 , n10591 , n10596 );
nor ( n10598 , n10585 , n10597 );
nand ( n10599 , n10579 , n10598 );
not ( n10600 , n10599 );
or ( n10601 , n2306 , n10600 );
or ( n10602 , n17 , n10217 );
nand ( n10603 , n10602 , n9406 );
and ( n10604 , n8044 , n10603 );
nor ( n10605 , n10604 , n10117 );
or ( n10606 , n42 , n10605 );
not ( n10607 , n9088 );
nand ( n10608 , n10607 , n10187 , n10185 , n10196 );
and ( n10609 , n10140 , n10608 );
not ( n10610 , n17 );
not ( n10611 , n10610 );
not ( n10612 , n10206 );
or ( n10613 , n10611 , n10612 );
nand ( n10614 , n10613 , n9406 );
and ( n10615 , n3299 , n10614 );
nor ( n10616 , n10609 , n10615 );
nand ( n10617 , n10601 , n10606 , n10616 );
and ( n10618 , n92 , n10170 );
not ( n10619 , n10160 );
nor ( n10620 , n10619 , n15 , n26 , n10001 );
nor ( n10621 , n10618 , n10620 , n9680 );
or ( n10622 , n6679 , n10621 );
not ( n10623 , n10392 );
or ( n10624 , n9829 , n9578 , n10577 );
not ( n10625 , n10232 );
and ( n10626 , n9579 , n10625 );
and ( n10627 , n2347 , n9280 );
nor ( n10628 , n10626 , n10627 );
nand ( n10629 , n10624 , n10628 );
nand ( n10630 , n10623 , n10629 );
nand ( n10631 , n10622 , n10630 );
not ( n10632 , n10147 );
not ( n10633 , n92 );
or ( n10634 , n9835 , n10304 );
not ( n10635 , n9348 );
and ( n10636 , n10074 , n10635 );
nand ( n10637 , n551 , n9849 );
or ( n10638 , n9835 , n10294 );
nand ( n10639 , n10638 , n10302 );
nand ( n10640 , n10637 , n10639 );
nor ( n10641 , n10636 , n10640 );
nand ( n10642 , n10634 , n10641 );
not ( n10643 , n10642 );
or ( n10644 , n10633 , n10643 );
nand ( n10645 , n10644 , n9681 );
not ( n10646 , n10645 );
or ( n10647 , n10632 , n10646 );
nand ( n10648 , n10647 , n10114 );
nor ( n10649 , n10617 , n10631 , n10648 );
not ( n10650 , n9806 );
not ( n10651 , n9583 );
not ( n10652 , n10589 );
not ( n10653 , n9088 );
nand ( n10654 , n10652 , n10653 );
and ( n10655 , n15 , n10651 , n10654 );
nor ( n10656 , n10655 , n10629 );
and ( n10657 , n450 , n10599 );
not ( n10658 , n14 );
and ( n10659 , n10658 , n10603 );
nor ( n10660 , n10657 , n10659 );
nand ( n10661 , n10656 , n10660 );
and ( n10662 , n10650 , n10661 );
and ( n10663 , n10160 , n1382 , n10573 );
not ( n10664 , n10575 );
or ( n10665 , n10664 , n10166 );
nand ( n10666 , n10665 , n10181 );
nor ( n10667 , n10663 , n10666 );
and ( n10668 , n9432 , n10206 );
not ( n10669 , n32 );
and ( n10670 , n10669 , n9478 , n4346 );
nor ( n10671 , n10670 , n9327 );
nor ( n10672 , n10668 , n10671 );
and ( n10673 , n9428 , n10198 );
and ( n10674 , n234 , n9347 );
not ( n10675 , n10166 );
nor ( n10676 , n10674 , n10675 );
or ( n10677 , n32 , n10676 );
nand ( n10678 , n10677 , n10167 );
and ( n10679 , n10573 , n10678 );
nor ( n10680 , n10673 , n10679 );
nand ( n10681 , n10667 , n10672 , n10680 );
and ( n10682 , n10155 , n10681 );
nand ( n10683 , n32 , n10312 );
and ( n10684 , n10471 , n10683 );
not ( n10685 , n32 );
nand ( n10686 , n10685 , n10319 );
nand ( n10687 , n10684 , n10318 , n10686 );
and ( n10688 , n9974 , n10687 );
nor ( n10689 , n10662 , n10682 , n10688 );
not ( n10690 , n9898 );
and ( n10691 , n9428 , n10687 );
or ( n10692 , n32 , n10288 );
not ( n10693 , n10247 );
not ( n10694 , n10282 );
or ( n10695 , n10693 , n10694 );
nand ( n10696 , n10695 , n10431 );
nand ( n10697 , n10692 , n10696 );
nor ( n10698 , n10697 , n10642 );
or ( n10699 , n9313 , n10698 );
nand ( n10700 , n10699 , n10322 );
or ( n10701 , n35 , n9917 );
not ( n10702 , n32 );
nand ( n10703 , n10701 , n10702 );
nand ( n10704 , n22 , n10703 );
nand ( n10705 , n10074 , n4374 );
and ( n10706 , n10704 , n10705 );
nor ( n10707 , n10706 , n9483 );
nor ( n10708 , n10691 , n10700 , n10707 );
not ( n10709 , n10708 );
and ( n10710 , n10690 , n10709 );
not ( n10711 , n17 );
not ( n10712 , n10711 );
not ( n10713 , n10697 );
or ( n10714 , n10712 , n10713 );
nand ( n10715 , n10714 , n9406 );
and ( n10716 , n6835 , n10715 );
nor ( n10717 , n10710 , n10716 );
not ( n10718 , n10028 );
or ( n10719 , n9484 , n9566 );
not ( n10720 , n9762 );
or ( n10721 , n9484 , n10720 );
nand ( n10722 , n10721 , n10001 );
not ( n10723 , n10358 );
and ( n10724 , n10722 , n10723 );
not ( n10725 , n10001 );
not ( n10726 , n10361 );
or ( n10727 , n10725 , n10726 );
not ( n10728 , n9844 );
nand ( n10729 , n10723 , n255 , n10728 );
nand ( n10730 , n10727 , n10729 );
nor ( n10731 , n10724 , n10730 );
nand ( n10732 , n10719 , n10731 , n10637 );
and ( n10733 , n9579 , n10732 );
not ( n10734 , n14 );
not ( n10735 , n32 );
and ( n10736 , n10735 , n10353 );
and ( n10737 , n10247 , n10347 );
nor ( n10738 , n10737 , n10430 );
nor ( n10739 , n10736 , n10738 );
or ( n10740 , n17 , n10739 );
nand ( n10741 , n10740 , n9406 );
and ( n10742 , n10734 , n10741 );
nor ( n10743 , n10733 , n10742 );
nand ( n10744 , n10074 , n10509 );
and ( n10745 , n10704 , n10744 );
nor ( n10746 , n10745 , n9483 );
not ( n10747 , n10746 );
nand ( n10748 , n10747 , n10341 );
or ( n10749 , n9313 , n10739 );
nand ( n10750 , n9432 , n10732 );
nand ( n10751 , n32 , n10330 );
and ( n10752 , n10471 , n10751 );
not ( n10753 , n32 );
nand ( n10754 , n10753 , n10337 );
nand ( n10755 , n10752 , n10336 , n10754 );
nand ( n10756 , n9428 , n10755 );
nand ( n10757 , n10749 , n10750 , n10756 );
or ( n10758 , n10748 , n10757 );
nand ( n10759 , n10758 , n450 );
nand ( n10760 , n10743 , n9585 , n10759 );
and ( n10761 , n10465 , n10336 );
nand ( n10762 , n10761 , n10751 , n10754 );
not ( n10763 , n10762 );
and ( n10764 , n10341 , n10749 );
nor ( n10765 , n10746 , n10741 );
and ( n10766 , n10764 , n10765 , n9500 , n10750 );
nand ( n10767 , n10763 , n10766 , n10756 );
nand ( n10768 , n10760 , n10767 );
not ( n10769 , n10768 );
and ( n10770 , n10718 , n10769 );
and ( n10771 , n10384 , n10760 );
nor ( n10772 , n10770 , n10771 );
nand ( n10773 , n10649 , n10689 , n10717 , n10772 );
nand ( n10774 , n10571 , n10773 );
nand ( n10775 , n10494 , n10569 , n10570 , n10774 );
and ( n10776 , n10424 , n10775 );
not ( n10777 , n18 );
not ( n10778 , n10777 );
nand ( n10779 , n10518 , n9709 );
or ( n10780 , n35 , n9738 );
nand ( n10781 , n10780 , n32 );
not ( n10782 , n10781 );
not ( n10783 , n9742 );
or ( n10784 , n10782 , n10783 );
or ( n10785 , n7369 , n9721 );
nand ( n10786 , n10785 , n10431 );
nand ( n10787 , n10784 , n10786 );
nand ( n10788 , n9432 , n10787 );
nand ( n10789 , n32 , n9696 );
and ( n10790 , n10471 , n10789 );
not ( n10791 , n32 );
nand ( n10792 , n10791 , n9705 );
nand ( n10793 , n10790 , n9704 , n10792 );
nand ( n10794 , n9428 , n10793 );
not ( n10795 , n9484 );
not ( n10796 , n9764 );
or ( n10797 , n10795 , n10796 );
nand ( n10798 , n10797 , n9835 );
not ( n10799 , n10798 );
not ( n10800 , n9772 );
or ( n10801 , n10799 , n10800 );
nand ( n10802 , n7370 , n9365 );
not ( n10803 , n9759 );
or ( n10804 , n10802 , n10803 );
nand ( n10805 , n10804 , n9835 );
nand ( n10806 , n10801 , n10805 );
nand ( n10807 , n9432 , n10806 );
nand ( n10808 , n10788 , n10794 , n10807 );
nor ( n10809 , n10779 , n10808 );
or ( n10810 , n2065 , n10809 );
and ( n10811 , n9579 , n10806 );
not ( n10812 , n17 );
and ( n10813 , n10812 , n10787 );
nor ( n10814 , n10813 , n9284 );
or ( n10815 , n14 , n10814 );
nand ( n10816 , n10815 , n9585 );
nor ( n10817 , n10811 , n10816 );
nand ( n10818 , n10810 , n10817 );
not ( n10819 , n10818 );
or ( n10820 , n10819 , n2384 , n2955 );
not ( n10821 , n17 );
or ( n10822 , n9637 , n32 );
not ( n10823 , n9617 );
or ( n10824 , n10430 , n10823 );
nand ( n10825 , n22 , n9621 );
not ( n10826 , n35 );
and ( n10827 , n10825 , n10826 , n9635 );
nor ( n10828 , n10430 , n118 );
nor ( n10829 , n10827 , n10828 );
nand ( n10830 , n10822 , n10824 , n10829 );
and ( n10831 , n10821 , n10830 );
nor ( n10832 , n10831 , n9284 );
or ( n10833 , n6368 , n10832 );
nand ( n10834 , n10820 , n10833 );
and ( n10835 , n20 , n10118 );
and ( n10836 , n2066 , n9445 );
nand ( n10837 , n20 , n9686 );
nand ( n10838 , n32 , n9598 );
and ( n10839 , n10471 , n10838 );
not ( n10840 , n32 );
nand ( n10841 , n10840 , n9606 );
and ( n10842 , n10839 , n9605 , n10841 );
or ( n10843 , n10837 , n2384 , n10842 );
not ( n10844 , n9445 );
or ( n10845 , n3089 , n10844 );
nand ( n10846 , n10843 , n10845 );
nor ( n10847 , n10835 , n10836 , n10846 );
and ( n10848 , n9978 , n10671 );
not ( n10849 , n9984 );
or ( n10850 , n10849 , n9994 );
and ( n10851 , n10128 , n10132 );
or ( n10852 , n10123 , n10851 );
or ( n10853 , n9983 , n10013 );
nand ( n10854 , n10850 , n10852 , n10853 );
nor ( n10855 , n10848 , n10854 );
or ( n10856 , n9999 , n10013 );
nand ( n10857 , n10855 , n10024 , n10021 , n10856 );
and ( n10858 , n20 , n10857 );
not ( n10859 , n9250 );
and ( n10860 , n10427 , n10859 );
not ( n10861 , n9238 );
nand ( n10862 , n10247 , n10861 );
and ( n10863 , n10431 , n10862 );
nor ( n10864 , n10860 , n10863 );
or ( n10865 , n17 , n10864 );
and ( n10866 , n10001 , n9273 );
and ( n10867 , n9835 , n10439 );
nor ( n10868 , n10866 , n10867 );
or ( n10869 , n692 , n10868 );
nand ( n10870 , n10865 , n10869 , n9285 );
and ( n10871 , n1919 , n10870 );
or ( n10872 , n21 , n1939 , n10851 );
or ( n10873 , n21 , n963 , n9290 );
nand ( n10874 , n10872 , n10873 );
nor ( n10875 , n10858 , n10871 , n10874 );
not ( n10876 , n9964 );
and ( n10877 , n10001 , n10876 );
nand ( n10878 , n7370 , n9942 );
not ( n10879 , n9958 );
or ( n10880 , n10878 , n10879 );
nand ( n10881 , n10880 , n9835 );
not ( n10882 , n9963 );
nand ( n10883 , n10881 , n10882 );
nor ( n10884 , n10877 , n10883 );
or ( n10885 , n15 , n10884 );
nand ( n10886 , n10885 , n9683 );
and ( n10887 , n10886 , n2245 , n2066 );
not ( n10888 , n10837 );
not ( n10889 , n32 );
or ( n10890 , n10889 , n9903 );
not ( n10891 , n32 );
nand ( n10892 , n10891 , n9912 );
nand ( n10893 , n10471 , n10890 , n9911 , n10892 );
and ( n10894 , n2816 , n10888 , n10893 );
nor ( n10895 , n10887 , n10894 );
not ( n10896 , n17 );
not ( n10897 , n10896 );
or ( n10898 , n9935 , n32 );
or ( n10899 , n10430 , n9924 );
nand ( n10900 , n22 , n9933 );
and ( n10901 , n10900 , n35 , n9929 );
nor ( n10902 , n10901 , n10828 );
nand ( n10903 , n10898 , n10899 , n10902 );
not ( n10904 , n10903 );
or ( n10905 , n10897 , n10904 );
nand ( n10906 , n10905 , n9406 );
and ( n10907 , n2389 , n10906 );
and ( n10908 , n9484 , n9664 );
nor ( n10909 , n10908 , n10001 );
or ( n10910 , n10909 , n9669 );
not ( n10911 , n9658 );
nor ( n10912 , n10911 , n10802 );
or ( n10913 , n10001 , n10912 );
nand ( n10914 , n10910 , n10913 );
and ( n10915 , n92 , n10914 );
nor ( n10916 , n10915 , n9682 );
nor ( n10917 , n10916 , n2244 , n3089 );
nor ( n10918 , n10907 , n10917 );
nand ( n10919 , n10847 , n10875 , n10895 , n10918 );
nor ( n10920 , n10834 , n10919 );
not ( n10921 , n10789 );
nor ( n10922 , n1387 , n10921 );
nand ( n10923 , n10922 , n9704 , n10792 );
not ( n10924 , n10923 );
or ( n10925 , n10924 , n10817 );
not ( n10926 , n2065 );
not ( n10927 , n10817 );
or ( n10928 , n10926 , n10927 );
not ( n10929 , n10809 );
nand ( n10930 , n10928 , n10929 );
not ( n10931 , n9500 );
not ( n10932 , n10814 );
or ( n10933 , n10931 , n10932 );
nand ( n10934 , n10933 , n10818 );
nand ( n10935 , n10925 , n10930 , n10934 );
and ( n10936 , n10935 , n2487 , n2385 );
not ( n10937 , n10842 );
nand ( n10938 , n10937 , n9428 );
or ( n10939 , n10830 , n10914 );
nand ( n10940 , n10939 , n9432 );
nand ( n10941 , n9609 , n10559 , n10938 , n10940 );
and ( n10942 , n10941 , n2229 , n3090 );
nor ( n10943 , n10936 , n10942 );
not ( n10944 , n2629 );
and ( n10945 , n9428 , n10893 );
nor ( n10946 , n10945 , n10707 );
not ( n10947 , n9914 );
not ( n10948 , n10884 );
or ( n10949 , n10903 , n10948 );
nand ( n10950 , n10949 , n9432 );
and ( n10951 , n10946 , n10947 , n10950 );
not ( n10952 , n10951 );
and ( n10953 , n10944 , n10952 );
nand ( n10954 , n7370 , n9323 );
and ( n10955 , n32 , n10954 );
not ( n10956 , n32 );
and ( n10957 , n10956 , n9307 );
nor ( n10958 , n10955 , n10957 );
or ( n10959 , n21 , n10958 );
not ( n10960 , n10958 );
and ( n10961 , n9428 , n10960 );
and ( n10962 , n10864 , n10868 );
nor ( n10963 , n10962 , n9313 );
nand ( n10964 , n10478 , n9331 );
nor ( n10965 , n10961 , n10963 , n10964 );
nand ( n10966 , n10959 , n10965 );
and ( n10967 , n942 , n10966 );
nor ( n10968 , n10953 , n10967 );
not ( n10969 , n16 );
not ( n10970 , n2487 );
nor ( n10971 , n10970 , n19 );
not ( n10972 , n14 );
not ( n10973 , n17 );
not ( n10974 , n10973 );
not ( n10975 , n9818 );
not ( n10976 , n10975 );
or ( n10977 , n10974 , n10976 );
nand ( n10978 , n10977 , n9406 );
and ( n10979 , n10972 , n10978 );
or ( n10980 , n9578 , n9851 );
nand ( n10981 , n10980 , n9585 );
nor ( n10982 , n10979 , n10981 );
or ( n10983 , n9500 , n10982 );
not ( n10984 , n2065 );
not ( n10985 , n10982 );
or ( n10986 , n10984 , n10985 );
nor ( n10987 , n9866 , n9876 );
not ( n10988 , n10987 );
and ( n10989 , n9428 , n10988 );
and ( n10990 , n9432 , n10975 );
nor ( n10991 , n10989 , n10990 );
or ( n10992 , n9313 , n9851 );
nand ( n10993 , n10992 , n9881 );
nor ( n10994 , n10583 , n10993 );
nand ( n10995 , n10991 , n10994 );
nand ( n10996 , n10986 , n10995 );
or ( n10997 , n10978 , n10988 );
not ( n10998 , n450 );
not ( n10999 , n10995 );
or ( n11000 , n10998 , n10999 );
nand ( n11001 , n11000 , n10982 );
nand ( n11002 , n10997 , n11001 );
nand ( n11003 , n10983 , n10996 , n11002 );
nand ( n11004 , n10969 , n10971 , n11003 );
and ( n11005 , n10001 , n10087 );
not ( n11006 , n10081 );
or ( n11007 , n10878 , n11006 );
nand ( n11008 , n11007 , n9835 );
nand ( n11009 , n11008 , n10086 );
nor ( n11010 , n11005 , n11009 );
or ( n11011 , n9578 , n11010 );
not ( n11012 , n35 );
not ( n11013 , n10062 );
or ( n11014 , n11012 , n11013 );
nand ( n11015 , n11014 , n32 );
and ( n11016 , n11015 , n10065 );
not ( n11017 , n10060 );
and ( n11018 , n7370 , n11017 );
nor ( n11019 , n11018 , n10430 );
nor ( n11020 , n11016 , n11019 );
not ( n11021 , n11020 );
not ( n11022 , n17 );
and ( n11023 , n11021 , n11022 );
nor ( n11024 , n11023 , n9284 );
or ( n11025 , n14 , n11024 );
nand ( n11026 , n11011 , n11025 , n9585 );
not ( n11027 , n11026 );
nand ( n11028 , n32 , n10031 );
not ( n11029 , n32 );
nand ( n11030 , n11029 , n10042 );
nand ( n11031 , n10471 , n11028 , n10041 , n11030 );
nand ( n11032 , n9428 , n11031 );
not ( n11033 , n11032 );
not ( n11034 , n10032 );
or ( n11035 , n10746 , n11034 );
and ( n11036 , n11020 , n11010 );
nor ( n11037 , n11036 , n9313 );
nor ( n11038 , n11035 , n11037 );
not ( n11039 , n11038 );
or ( n11040 , n11033 , n11039 );
nand ( n11041 , n11040 , n450 );
nand ( n11042 , n11027 , n11041 );
not ( n11043 , n11042 );
or ( n11044 , n2815 , n11043 );
not ( n11045 , n11001 );
or ( n11046 , n1407 , n11045 );
nand ( n11047 , n11044 , n11046 );
nand ( n11048 , n2954 , n11047 );
and ( n11049 , n10465 , n11028 );
nand ( n11050 , n11049 , n10041 , n11030 );
nand ( n11051 , n11050 , n11026 );
or ( n11052 , n11026 , n450 );
not ( n11053 , n9428 );
not ( n11054 , n11050 );
or ( n11055 , n11053 , n11054 );
nand ( n11056 , n11055 , n11038 );
nand ( n11057 , n11052 , n11056 );
not ( n11058 , n9500 );
not ( n11059 , n11024 );
or ( n11060 , n11058 , n11059 );
nand ( n11061 , n11060 , n11042 );
and ( n11062 , n11051 , n11057 , n11061 );
not ( n11063 , n11062 );
nand ( n11064 , n16 , n10971 , n11063 );
and ( n11065 , n11004 , n11048 , n11064 );
nand ( n11066 , n10920 , n10943 , n10968 , n11065 );
not ( n11067 , n11066 );
or ( n11068 , n10778 , n11067 );
nand ( n11069 , n9470 , n9686 , n9442 );
nand ( n11070 , n11068 , n11069 );
nor ( n11071 , n10776 , n11070 );
nand ( n11072 , n9448 , n9804 , n10423 , n11071 );
and ( n11073 , n2510 , n11072 );
or ( n11074 , n1888 , n9672 );
nor ( n11075 , n2244 , n2384 );
not ( n11076 , n11075 );
not ( n11077 , n9684 );
or ( n11078 , n11076 , n11077 );
nand ( n11079 , n11074 , n11078 );
and ( n11080 , n1582 , n11079 );
and ( n11081 , n96 , n9968 );
and ( n11082 , n2235 , n10136 );
nor ( n11083 , n11081 , n11082 );
or ( n11084 , n11083 , n1599 );
not ( n11085 , n14 );
nor ( n11086 , n11085 , n2384 );
and ( n11087 , n11086 , n9676 );
and ( n11088 , n1373 , n9338 );
nor ( n11089 , n11087 , n11088 );
or ( n11090 , n1984 , n11089 );
nand ( n11091 , n6674 , n3425 );
not ( n11092 , n10149 );
or ( n11093 , n11091 , n11092 );
nand ( n11094 , n11084 , n11090 , n11093 );
nor ( n11095 , n11080 , n11094 );
nor ( n11096 , n21 , n295 );
and ( n11097 , n9976 , n3425 , n11096 );
not ( n11098 , n21 );
not ( n11099 , n9088 );
not ( n11100 , n11099 );
not ( n11101 , n11100 );
nand ( n11102 , n11101 , n10133 );
and ( n11103 , n11098 , n2003 , n11102 );
nor ( n11104 , n11097 , n11103 );
or ( n11105 , n10134 , n10025 );
nand ( n11106 , n11105 , n1582 );
nand ( n11107 , n11095 , n11104 , n11106 );
or ( n11108 , n16 , n2862 , n9896 );
or ( n11109 , n2864 , n10107 );
nand ( n11110 , n11108 , n11109 );
not ( n11111 , n11110 );
nor ( n11112 , n1984 , n1375 );
and ( n11113 , n11112 , n9334 );
and ( n11114 , n2228 , n970 );
not ( n11115 , n19 );
nor ( n11116 , n11114 , n11115 , n21 );
not ( n11117 , n11116 );
not ( n11118 , n11101 );
buf ( n11119 , n11118 );
not ( n11120 , n11119 );
or ( n11121 , n11117 , n1984 , n11120 );
not ( n11122 , n4323 );
nand ( n11123 , n11122 , n11096 );
or ( n11124 , n1599 , n11123 );
nand ( n11125 , n11121 , n11124 );
nor ( n11126 , n1984 , n1888 , n21 , n9607 );
nor ( n11127 , n11113 , n11125 , n11126 );
and ( n11128 , n5121 , n9440 );
nor ( n11129 , n21 , n591 );
and ( n11130 , n11129 , n9470 );
nor ( n11131 , n11128 , n11130 );
not ( n11132 , n11123 );
and ( n11133 , n453 , n11132 );
not ( n11134 , n20 );
nand ( n11135 , n11134 , n11116 );
nor ( n11136 , n10653 , n11135 );
nor ( n11137 , n11133 , n11136 );
nand ( n11138 , n2243 , n10401 );
and ( n11139 , n11131 , n11137 , n11138 );
and ( n11140 , n453 , n11096 );
and ( n11141 , n11140 , n10406 );
and ( n11142 , n6676 , n10398 );
nor ( n11143 , n11141 , n11142 );
not ( n11144 , n20 );
not ( n11145 , n1373 );
not ( n11146 , n9286 );
or ( n11147 , n11145 , n11146 );
nand ( n11148 , n11086 , n9407 );
nand ( n11149 , n11147 , n11148 );
nand ( n11150 , n11144 , n11149 );
nand ( n11151 , n11075 , n9373 );
nand ( n11152 , n764 , n9493 );
and ( n11153 , n11151 , n11152 );
nor ( n11154 , n11153 , n20 );
not ( n11155 , n11154 );
and ( n11156 , n11139 , n11143 , n11150 , n11155 );
nor ( n11157 , n2244 , n1931 );
and ( n11158 , n11157 , n10412 );
and ( n11159 , n3146 , n10418 );
nor ( n11160 , n11158 , n11159 );
nand ( n11161 , n8976 , n10212 );
and ( n11162 , n11156 , n11160 , n11161 );
not ( n11163 , n9588 );
or ( n11164 , n1931 , n10274 );
and ( n11165 , n1547 , n10117 );
not ( n11166 , n4323 );
not ( n11167 , n11166 );
nand ( n11168 , n11167 , n10188 , n10189 , n10199 );
nand ( n11169 , n11165 , n11168 );
nand ( n11170 , n11164 , n11169 );
or ( n11171 , n2186 , n10378 );
nor ( n11172 , n6286 , n10324 );
not ( n11173 , n11172 );
nand ( n11174 , n11171 , n11173 );
nor ( n11175 , n11170 , n11174 );
nand ( n11176 , n11162 , n11163 , n11175 );
and ( n11177 , n18 , n11176 );
and ( n11178 , n9591 , n9793 );
nor ( n11179 , n11177 , n11178 );
nand ( n11180 , n11111 , n11127 , n11179 );
nor ( n11181 , n11107 , n11180 );
nand ( n11182 , n1406 , n10857 );
nor ( n11183 , n6675 , n1315 );
and ( n11184 , n11183 , n10886 );
nor ( n11185 , n3471 , n1375 );
and ( n11186 , n11185 , n10966 );
nor ( n11187 , n11184 , n11186 );
and ( n11188 , n11182 , n11187 );
not ( n11189 , n11120 );
not ( n11190 , n11189 );
nand ( n11191 , n1406 , n11116 );
or ( n11192 , n11190 , n11191 );
not ( n11193 , n21 );
and ( n11194 , n11193 , n11189 , n1319 );
nand ( n11195 , n10653 , n10851 );
not ( n11196 , n11195 );
not ( n11197 , n14 );
nor ( n11198 , n11196 , n11197 , n21 , n8717 );
nor ( n11199 , n11194 , n11198 );
not ( n11200 , n16 );
and ( n11201 , n11200 , n6761 , n11003 );
nor ( n11202 , n3460 , n10951 );
nor ( n11203 , n11201 , n11202 );
and ( n11204 , n11188 , n11192 , n11199 , n11203 );
not ( n11205 , n2235 );
not ( n11206 , n10906 );
or ( n11207 , n11205 , n11206 );
nand ( n11208 , n11096 , n10893 );
nand ( n11209 , n11207 , n11208 );
and ( n11210 , n1314 , n11209 );
not ( n11211 , n1406 );
nor ( n11212 , n11211 , n1888 , n10842 , n21 );
not ( n11213 , n10832 );
and ( n11214 , n11086 , n11213 );
and ( n11215 , n1373 , n10870 );
nor ( n11216 , n11214 , n11215 );
nor ( n11217 , n3471 , n11216 );
nor ( n11218 , n11210 , n11212 , n11217 );
nor ( n11219 , n6762 , n11062 );
not ( n11220 , n764 );
not ( n11221 , n10941 );
or ( n11222 , n11220 , n11221 );
or ( n11223 , n11076 , n10916 );
nand ( n11224 , n11222 , n11223 );
nand ( n11225 , n1406 , n11224 );
nand ( n11226 , n8631 , n10935 );
and ( n11227 , n11165 , n10608 );
nand ( n11228 , n2243 , n10715 );
nand ( n11229 , n11137 , n11228 );
nor ( n11230 , n11227 , n11229 );
and ( n11231 , n5121 , n10481 );
and ( n11232 , n11129 , n10498 );
nor ( n11233 , n11231 , n11232 );
and ( n11234 , n1373 , n10446 );
and ( n11235 , n11086 , n10491 );
nor ( n11236 , n11234 , n11235 );
nor ( n11237 , n20 , n11236 );
not ( n11238 , n11237 );
and ( n11239 , n8976 , n10681 );
not ( n11240 , n3146 );
not ( n11241 , n10614 );
or ( n11242 , n11240 , n11241 );
not ( n11243 , n11157 );
or ( n11244 , n11243 , n10621 );
nand ( n11245 , n11242 , n11244 );
nor ( n11246 , n11239 , n11245 );
nand ( n11247 , n11230 , n11233 , n11238 , n11246 );
and ( n11248 , n3256 , n10661 );
and ( n11249 , n11140 , n10687 );
nor ( n11250 , n11248 , n11249 );
or ( n11251 , n6286 , n10708 );
nand ( n11252 , n11075 , n10459 );
nand ( n11253 , n764 , n10566 );
and ( n11254 , n11252 , n11253 );
nor ( n11255 , n11254 , n20 );
not ( n11256 , n11255 );
and ( n11257 , n11250 , n11251 , n11256 );
not ( n11258 , n2186 );
not ( n11259 , n10768 );
and ( n11260 , n11258 , n11259 );
and ( n11261 , n6676 , n10645 );
nor ( n11262 , n11260 , n11261 );
nand ( n11263 , n2458 , n10553 );
nand ( n11264 , n11257 , n11262 , n11263 );
or ( n11265 , n11247 , n11264 );
not ( n11266 , n18 );
nand ( n11267 , n11265 , n11266 );
nand ( n11268 , n11225 , n11226 , n11267 );
nor ( n11269 , n11219 , n11268 );
nand ( n11270 , n11181 , n11204 , n11218 , n11269 );
not ( n11271 , n11270 );
nor ( n11272 , n2731 , n11271 );
nor ( n11273 , n11073 , n11272 );
nand ( n11274 , n1582 , n3747 );
not ( n11275 , n11274 );
not ( n11276 , n10134 );
not ( n11277 , n10025 );
nand ( n11278 , n11276 , n11089 , n11277 , n10150 );
and ( n11279 , n11275 , n11278 );
not ( n11280 , n11116 );
not ( n11281 , n11079 );
and ( n11282 , n11280 , n11281 );
nor ( n11283 , n11282 , n11274 );
and ( n11284 , n3748 , n9591 , n9795 );
nor ( n11285 , n11279 , n11283 , n11284 );
not ( n11286 , n18 );
not ( n11287 , n3748 );
nor ( n11288 , n11286 , n11287 );
or ( n11289 , n1931 , n10393 );
not ( n11290 , n2261 );
nand ( n11291 , n11290 , n10398 );
not ( n11292 , n9973 );
not ( n11293 , n11117 );
or ( n11294 , n11292 , n11293 );
not ( n11295 , n20 );
nand ( n11296 , n11294 , n11295 );
and ( n11297 , n11291 , n11296 , n11150 );
nand ( n11298 , n11289 , n11297 );
not ( n11299 , n11298 );
and ( n11300 , n454 , n10375 );
nor ( n11301 , n11300 , n11172 , n11154 );
not ( n11302 , n9439 );
nand ( n11303 , n5121 , n11302 );
and ( n11304 , n11301 , n11303 , n11138 , n9587 );
nand ( n11305 , n11299 , n11304 , n11160 , n11161 );
and ( n11306 , n11288 , n11305 );
not ( n11307 , n10112 );
and ( n11308 , n11275 , n11307 );
nor ( n11309 , n11306 , n11308 );
nand ( n11310 , n9968 , n3748 , n3686 );
not ( n11311 , n10965 );
and ( n11312 , n11185 , n11311 );
nand ( n11313 , n11191 , n11182 );
nor ( n11314 , n11312 , n11313 );
not ( n11315 , n18 );
not ( n11316 , n20 );
nor ( n11317 , n11316 , n6834 );
nand ( n11318 , n11315 , n11317 , n10906 );
and ( n11319 , n10886 , n1406 , n10147 );
nor ( n11320 , n11319 , n11217 );
nand ( n11321 , n11314 , n11318 , n11320 );
and ( n11322 , n8631 , n10818 );
or ( n11323 , n1913 , n10951 );
nand ( n11324 , n11323 , n11225 );
nor ( n11325 , n11322 , n11324 );
not ( n11326 , n18 );
nand ( n11327 , n11326 , n2438 , n9686 );
nand ( n11328 , n1406 , n11047 );
not ( n11329 , n18 );
and ( n11330 , n8125 , n10599 );
not ( n11331 , n10645 );
or ( n11332 , n2261 , n11331 );
nand ( n11333 , n11332 , n11135 , n11228 );
and ( n11334 , n9973 , n10605 );
nor ( n11335 , n11334 , n20 );
nor ( n11336 , n11330 , n11333 , n11335 );
not ( n11337 , n10480 );
and ( n11338 , n5121 , n11337 );
and ( n11339 , n3256 , n10629 );
nor ( n11340 , n11338 , n11339 );
and ( n11341 , n11340 , n11246 , n11251 );
nor ( n11342 , n11237 , n11255 );
and ( n11343 , n454 , n10760 );
and ( n11344 , n2458 , n10544 );
nor ( n11345 , n11343 , n11344 );
nand ( n11346 , n11336 , n11341 , n11342 , n11345 );
nand ( n11347 , n11329 , n11346 );
nand ( n11348 , n11325 , n11327 , n11328 , n11347 );
or ( n11349 , n11321 , n11348 );
nand ( n11350 , n11349 , n3748 );
and ( n11351 , n11309 , n11310 , n11350 );
and ( n11352 , n3748 , n3425 , n9686 );
or ( n11353 , n9333 , n1375 , n11274 );
or ( n11354 , n11274 , n10137 );
nand ( n11355 , n11353 , n11354 );
nor ( n11356 , n11352 , n11355 );
not ( n11357 , n3748 );
nand ( n11358 , n11357 , n11270 );
nand ( n11359 , n11285 , n11351 , n11356 , n11358 );
nand ( n11360 , n2299 , n3 , n11359 );
nand ( n11361 , n11273 , n4262 , n11360 );
not ( n11362 , n11359 );
not ( n11363 , n2300 );
not ( n11364 , n11358 );
not ( n11365 , n11364 );
or ( n11366 , n11363 , n11365 );
nand ( n11367 , n2889 , n1971 , n11072 );
nand ( n11368 , n11366 , n11367 );
not ( n11369 , n11368 );
nand ( n11370 , n11362 , n11369 );
or ( n11371 , n11361 , n11370 );
not ( n11372 , n21 );
not ( n11373 , n11372 );
not ( n11374 , n4262 );
and ( n11375 , n11373 , n11374 );
nand ( n11376 , n4 , n4225 );
not ( n11377 , n11376 );
and ( n11378 , n11377 , n11362 );
nor ( n11379 , n11375 , n11378 );
not ( n11380 , n11273 );
nor ( n11381 , n11380 , n11368 );
nand ( n11382 , n11381 , n9012 , n11360 );
nand ( n11383 , n11371 , n11379 , n11382 );
not ( n11384 , n3748 );
nand ( n11385 , n4249 , n11384 );
nor ( n11386 , n18 , n4240 , n11385 );
not ( n11387 , n20 );
not ( n11388 , n21 );
nor ( n11389 , n11388 , n5061 );
nand ( n11390 , n11389 , n2123 );
nor ( n11391 , n11387 , n11390 );
not ( n11392 , n11167 );
or ( n11393 , n11392 , n10988 );
nand ( n11394 , n11393 , n7809 );
and ( n11395 , n11391 , n11394 );
not ( n11396 , n448 );
and ( n11397 , n11396 , n11389 );
not ( n11398 , n11397 );
nor ( n11399 , n2391 , n11398 );
not ( n11400 , n11399 );
nand ( n11401 , n7809 , n11195 );
not ( n11402 , n11401 );
or ( n11403 , n11400 , n11402 );
nand ( n11404 , n11389 , n942 );
not ( n11405 , n10653 );
not ( n11406 , n10958 );
or ( n11407 , n11405 , n11406 );
nand ( n11408 , n11407 , n7809 );
not ( n11409 , n11408 );
or ( n11410 , n11404 , n11409 );
nand ( n11411 , n11403 , n11410 );
or ( n11412 , n7809 , n21 );
or ( n11413 , n998 , n11412 );
not ( n11414 , n21 );
not ( n11415 , n11414 );
not ( n11416 , n8616 );
or ( n11417 , n11415 , n11416 );
not ( n11418 , n21 );
nand ( n11419 , n11418 , n7809 );
nand ( n11420 , n11417 , n11419 );
and ( n11421 , n11420 , n11401 );
not ( n11422 , n21 );
nor ( n11423 , n7809 , n10851 );
and ( n11424 , n11422 , n11423 );
nor ( n11425 , n11421 , n11424 );
and ( n11426 , n11413 , n11425 );
not ( n11427 , n2781 );
nand ( n11428 , n20 , n11427 );
not ( n11429 , n3299 );
or ( n11430 , n11428 , n11429 );
nor ( n11431 , n11426 , n11430 );
nor ( n11432 , n11395 , n11411 , n11431 );
nor ( n11433 , n6368 , n11398 );
not ( n11434 , n11433 );
not ( n11435 , n11392 );
not ( n11436 , n11435 );
not ( n11437 , n10838 );
not ( n11438 , n9605 );
not ( n11439 , n10841 );
nor ( n11440 , n11437 , n1387 , n11438 , n11439 );
not ( n11441 , n11440 );
or ( n11442 , n11436 , n11441 );
nand ( n11443 , n11442 , n7809 );
not ( n11444 , n11443 );
or ( n11445 , n11434 , n11444 );
nand ( n11446 , n2389 , n11397 );
nor ( n11447 , n1387 , n11100 );
nand ( n11448 , n11447 , n9911 , n10890 , n10892 );
nand ( n11449 , n7809 , n11448 );
not ( n11450 , n11449 );
or ( n11451 , n11446 , n11450 );
nand ( n11452 , n11445 , n11451 );
and ( n11453 , n11420 , n11394 );
not ( n11454 , n21 );
nor ( n11455 , n7809 , n10987 );
and ( n11456 , n11454 , n11455 );
nor ( n11457 , n11453 , n11456 );
and ( n11458 , n11413 , n11457 );
nor ( n11459 , n11458 , n8567 );
not ( n11460 , n21 );
nand ( n11461 , n43 , n10893 );
not ( n11462 , n11461 );
and ( n11463 , n11460 , n11462 );
and ( n11464 , n11420 , n11449 );
nor ( n11465 , n11463 , n11464 );
and ( n11466 , n11413 , n11465 );
or ( n11467 , n11428 , n6834 );
nor ( n11468 , n11466 , n11467 );
nor ( n11469 , n11452 , n11459 , n11468 );
nor ( n11470 , n3516 , n6368 );
not ( n11471 , n21 );
not ( n11472 , n11471 );
nor ( n11473 , n7809 , n10842 );
not ( n11474 , n11473 );
or ( n11475 , n11472 , n11474 );
and ( n11476 , n11420 , n11443 );
not ( n11477 , n11413 );
nor ( n11478 , n11476 , n11477 );
nand ( n11479 , n11475 , n11478 );
and ( n11480 , n11470 , n11479 );
and ( n11481 , n2530 , n11455 );
nor ( n11482 , n7809 , n17 );
not ( n11483 , n11482 );
nand ( n11484 , n20 , n11483 );
nand ( n11485 , n3299 , n11423 );
nor ( n11486 , n11484 , n11485 );
nor ( n11487 , n11481 , n11486 );
and ( n11488 , n11408 , n1919 , n10960 );
not ( n11489 , n23 );
not ( n11490 , n9498 );
and ( n11491 , n11489 , n11490 );
nor ( n11492 , n11491 , n7809 );
not ( n11493 , n17 );
or ( n11494 , n11493 , n6360 );
nand ( n11495 , n11494 , n1920 );
and ( n11496 , n11492 , n11495 );
nand ( n11497 , n17 , n11492 );
not ( n11498 , n11497 );
and ( n11499 , n11498 , n6369 );
not ( n11500 , n8044 );
not ( n11501 , n11492 );
or ( n11502 , n11500 , n11501 );
not ( n11503 , n19 );
nand ( n11504 , n11503 , n11482 );
nand ( n11505 , n11502 , n11504 );
and ( n11506 , n20 , n11505 );
nor ( n11507 , n11496 , n11499 , n11506 );
not ( n11508 , n11507 );
nor ( n11509 , n11488 , n11508 );
not ( n11510 , n11420 );
nor ( n11511 , n963 , n11510 );
nand ( n11512 , n11511 , n11408 );
nor ( n11513 , n21 , n1418 );
and ( n11514 , n11408 , n11513 , n10960 );
and ( n11515 , n8572 , n11477 );
nor ( n11516 , n11515 , n11482 );
nor ( n11517 , n912 , n11516 );
nor ( n11518 , n11514 , n11517 );
nand ( n11519 , n11487 , n11509 , n11512 , n11518 );
not ( n11520 , n11473 );
or ( n11521 , n6368 , n11482 , n11520 );
or ( n11522 , n11484 , n6834 , n11461 );
nand ( n11523 , n11521 , n11522 );
nor ( n11524 , n11480 , n11519 , n11523 );
not ( n11525 , n2386 );
not ( n11526 , n11412 );
and ( n11527 , n11526 , n10923 );
not ( n11528 , n11420 );
or ( n11529 , n11118 , n10923 );
nand ( n11530 , n11529 , n7809 );
not ( n11531 , n11530 );
or ( n11532 , n11528 , n11531 );
nand ( n11533 , n11532 , n11413 );
nor ( n11534 , n11527 , n11533 );
or ( n11535 , n3493 , n11534 );
and ( n11536 , n11397 , n11530 );
nand ( n11537 , n17 , n43 );
not ( n11538 , n11537 );
and ( n11539 , n11538 , n10923 );
nor ( n11540 , n11536 , n11539 );
nand ( n11541 , n11535 , n11540 , n11497 );
and ( n11542 , n11525 , n11541 );
and ( n11543 , n11526 , n11050 );
nor ( n11544 , n11392 , n11050 );
or ( n11545 , n43 , n11544 );
not ( n11546 , n11545 );
or ( n11547 , n11510 , n11546 );
nand ( n11548 , n11547 , n11413 );
nor ( n11549 , n11543 , n11548 );
or ( n11550 , n3516 , n11549 );
and ( n11551 , n11397 , n11545 );
and ( n11552 , n11538 , n11050 );
nor ( n11553 , n11551 , n11552 );
nand ( n11554 , n11550 , n11553 , n11497 );
and ( n11555 , n2549 , n11554 );
nor ( n11556 , n11542 , n11555 );
nand ( n11557 , n11432 , n11469 , n11524 , n11556 );
and ( n11558 , n11386 , n11557 );
not ( n11559 , n18 );
nor ( n11560 , n11559 , n4240 , n11385 );
or ( n11561 , n11119 , n9606 );
nand ( n11562 , n11561 , n7809 );
and ( n11563 , n11433 , n11562 );
not ( n11564 , n3493 );
nand ( n11565 , n9089 , n9706 );
and ( n11566 , n7809 , n11565 );
or ( n11567 , n11510 , n11566 );
or ( n11568 , n11412 , n9708 );
nand ( n11569 , n11567 , n11568 , n11413 );
and ( n11570 , n11564 , n11569 );
or ( n11571 , n11398 , n11566 );
or ( n11572 , n11537 , n9708 );
nand ( n11573 , n11571 , n11572 );
nor ( n11574 , n11570 , n11573 , n11498 );
or ( n11575 , n2386 , n11574 );
not ( n11576 , n11404 );
or ( n11577 , n11118 , n9307 );
nand ( n11578 , n11577 , n7809 );
not ( n11579 , n11578 );
not ( n11580 , n11579 );
and ( n11581 , n11576 , n11580 );
nor ( n11582 , n7809 , n1920 );
and ( n11583 , n11582 , n9307 );
nor ( n11584 , n11581 , n11583 );
nand ( n11585 , n11575 , n11584 , n11507 );
not ( n11586 , n11419 );
not ( n11587 , n11102 );
and ( n11588 , n11586 , n11587 );
nand ( n11589 , n8622 , n10133 );
and ( n11590 , n11526 , n11589 );
nor ( n11591 , n11588 , n11590 );
and ( n11592 , n11413 , n11591 );
nor ( n11593 , n11592 , n11430 );
nor ( n11594 , n11563 , n11585 , n11593 );
not ( n11595 , n11594 );
not ( n11596 , n3493 );
not ( n11597 , n11166 );
not ( n11598 , n10042 );
and ( n11599 , n11597 , n11598 );
nor ( n11600 , n11599 , n43 );
or ( n11601 , n11419 , n11600 );
not ( n11602 , n8620 );
not ( n11603 , n11602 );
nor ( n11604 , n11603 , n10042 );
or ( n11605 , n11412 , n11604 );
nand ( n11606 , n11601 , n11605 , n11413 );
and ( n11607 , n11596 , n11606 );
and ( n11608 , n11538 , n10042 );
or ( n11609 , n11398 , n11600 );
nand ( n11610 , n11609 , n11497 );
nor ( n11611 , n11607 , n11608 , n11610 );
or ( n11612 , n2564 , n11611 );
not ( n11613 , n11413 );
and ( n11614 , n11420 , n11562 );
not ( n11615 , n21 );
nor ( n11616 , n7809 , n9607 );
and ( n11617 , n11615 , n11616 );
nor ( n11618 , n11614 , n11617 );
not ( n11619 , n11618 );
or ( n11620 , n11613 , n11619 );
nand ( n11621 , n11620 , n11470 );
nand ( n11622 , n11612 , n11621 );
not ( n11623 , n11118 );
and ( n11624 , n11623 , n9879 );
nor ( n11625 , n11624 , n43 );
not ( n11626 , n11625 );
and ( n11627 , n11420 , n11626 );
not ( n11628 , n21 );
nor ( n11629 , n7809 , n9879 );
and ( n11630 , n11628 , n11629 );
nor ( n11631 , n11627 , n11630 );
and ( n11632 , n11413 , n11631 );
nor ( n11633 , n11632 , n8567 );
or ( n11634 , n11119 , n9912 );
nand ( n11635 , n11634 , n7809 );
and ( n11636 , n11420 , n11635 );
not ( n11637 , n21 );
nor ( n11638 , n7809 , n9975 );
and ( n11639 , n11637 , n11638 );
nor ( n11640 , n11636 , n11639 );
and ( n11641 , n11413 , n11640 );
nor ( n11642 , n11641 , n11467 );
nor ( n11643 , n11595 , n11622 , n11633 , n11642 );
nand ( n11644 , n7809 , n11102 );
and ( n11645 , n11399 , n11644 );
or ( n11646 , n10133 , n11537 , n2391 );
nand ( n11647 , n11317 , n11483 , n11638 );
nand ( n11648 , n11646 , n11647 );
nand ( n11649 , n11513 , n9307 );
or ( n11650 , n7809 , n11649 );
and ( n11651 , n11511 , n11578 );
nor ( n11652 , n11651 , n11517 );
nand ( n11653 , n11650 , n11652 );
nor ( n11654 , n11645 , n11648 , n11653 );
and ( n11655 , n11391 , n11626 );
and ( n11656 , n2530 , n11629 );
nor ( n11657 , n11655 , n11656 );
and ( n11658 , n6426 , n11483 , n11616 );
not ( n11659 , n11635 );
nor ( n11660 , n11446 , n11659 );
nor ( n11661 , n11658 , n11660 );
nand ( n11662 , n11643 , n11654 , n11657 , n11661 );
and ( n11663 , n11560 , n11662 );
nor ( n11664 , n11558 , n11663 );
nand ( n11665 , n7 , n9014 );
not ( n11666 , n11665 );
or ( n11667 , n6 , n11666 );
nand ( n11668 , n11667 , n43 );
or ( n11669 , n9088 , n9421 );
nand ( n11670 , n11669 , n7809 );
nand ( n11671 , n7918 , n781 , n309 , n11670 );
not ( n11672 , n11671 );
nand ( n11673 , n2467 , n3128 );
and ( n11674 , n11673 , n18 , n11538 );
and ( n11675 , n43 , n18 , n3345 );
nor ( n11676 , n11674 , n11675 );
not ( n11677 , n1891 );
nand ( n11678 , n11677 , n7918 );
not ( n11679 , n11678 );
or ( n11680 , n11100 , n9470 );
nand ( n11681 , n11680 , n7809 );
nand ( n11682 , n11679 , n3251 , n18 , n11681 );
nand ( n11683 , n11676 , n11682 );
not ( n11684 , n21 );
nor ( n11685 , n7809 , n9543 );
and ( n11686 , n11684 , n11685 );
not ( n11687 , n11420 );
or ( n11688 , n11166 , n9542 );
nand ( n11689 , n11688 , n7809 );
not ( n11690 , n11689 );
or ( n11691 , n11687 , n11690 );
nand ( n11692 , n11691 , n11413 );
nor ( n11693 , n11686 , n11692 );
not ( n11694 , n3516 );
nand ( n11695 , n18 , n11694 );
nor ( n11696 , n11693 , n11695 , n3128 );
not ( n11697 , n21 );
nor ( n11698 , n7809 , n9471 );
and ( n11699 , n11697 , n11698 );
and ( n11700 , n11420 , n11681 );
nor ( n11701 , n11700 , n11477 );
not ( n11702 , n11701 );
nor ( n11703 , n11699 , n11702 );
or ( n11704 , n11703 , n11695 , n2467 );
nand ( n11705 , n11679 , n2515 );
not ( n11706 , n18 );
not ( n11707 , n11689 );
or ( n11708 , n11705 , n11706 , n11707 );
nand ( n11709 , n11704 , n11708 );
nor ( n11710 , n11672 , n11683 , n11696 , n11709 );
not ( n11711 , n11642 );
nor ( n11712 , n11678 , n2391 );
and ( n11713 , n11712 , n11644 );
nor ( n11714 , n7919 , n963 );
and ( n11715 , n11714 , n11578 );
nor ( n11716 , n6368 , n11678 );
not ( n11717 , n11716 );
not ( n11718 , n11562 );
or ( n11719 , n11717 , n11718 );
not ( n11720 , n11428 );
not ( n11721 , n6726 );
nand ( n11722 , n11720 , n11606 , n11721 );
nand ( n11723 , n11719 , n11722 );
nor ( n11724 , n11713 , n11715 , n11723 );
nand ( n11725 , n11679 , n2389 );
not ( n11726 , n11725 );
not ( n11727 , n11659 );
and ( n11728 , n11726 , n11727 );
nor ( n11729 , n3516 , n2386 );
and ( n11730 , n11729 , n11569 );
nor ( n11731 , n11728 , n11730 );
nand ( n11732 , n11711 , n11724 , n11731 , n11621 );
nand ( n11733 , n11679 , n2549 );
or ( n11734 , n11733 , n11600 );
nor ( n11735 , n11678 , n2386 );
not ( n11736 , n11735 );
or ( n11737 , n11736 , n11566 );
nor ( n11738 , n7919 , n795 );
nand ( n11739 , n20 , n11738 );
or ( n11740 , n11739 , n11625 );
nand ( n11741 , n11734 , n11737 , n11740 );
and ( n11742 , n11538 , n2549 );
nor ( n11743 , n6426 , n11525 );
or ( n11744 , n11537 , n11743 );
or ( n11745 , n11537 , n2393 );
not ( n11746 , n20 );
not ( n11747 , n11504 );
nor ( n11748 , n7809 , n14 , n1407 );
nor ( n11749 , n11747 , n11748 );
or ( n11750 , n11746 , n11749 );
nand ( n11751 , n11744 , n11745 , n11750 );
nor ( n11752 , n11742 , n11751 , n11582 );
not ( n11753 , n11752 );
or ( n11754 , n11753 , n11633 , n11653 , n11593 );
or ( n11755 , n11732 , n11741 , n11754 );
nand ( n11756 , n11755 , n18 );
not ( n11757 , n21 );
and ( n11758 , n10471 , n9540 );
and ( n11759 , n11758 , n10501 , n10503 );
nor ( n11760 , n11759 , n7809 );
and ( n11761 , n11757 , n11760 );
not ( n11762 , n11392 );
not ( n11763 , n10504 );
and ( n11764 , n11762 , n11763 );
nor ( n11765 , n11764 , n43 );
not ( n11766 , n11765 );
and ( n11767 , n11420 , n11766 );
nor ( n11768 , n11767 , n11477 );
not ( n11769 , n11768 );
nor ( n11770 , n11761 , n11769 );
or ( n11771 , n11770 , n3516 , n3128 );
not ( n11772 , n3516 );
not ( n11773 , n20 );
nand ( n11774 , n43 , n10755 );
or ( n11775 , n21 , n11774 );
or ( n11776 , n11119 , n10762 );
nand ( n11777 , n11776 , n7809 );
and ( n11778 , n11420 , n11777 );
nor ( n11779 , n11778 , n11477 );
nand ( n11780 , n11775 , n11779 );
nand ( n11781 , n11772 , n11721 , n11773 , n11780 );
nand ( n11782 , n11771 , n11781 );
not ( n11783 , n3493 );
nand ( n11784 , n11783 , n3251 );
not ( n11785 , n11784 );
not ( n11786 , n10564 );
or ( n11787 , n11412 , n11786 );
and ( n11788 , n11623 , n11786 );
nor ( n11789 , n11788 , n43 );
or ( n11790 , n11510 , n11789 );
nand ( n11791 , n11790 , n11413 );
not ( n11792 , n11791 );
nand ( n11793 , n11787 , n11792 );
nand ( n11794 , n11785 , n11793 );
not ( n11795 , n11789 );
and ( n11796 , n11795 , n11679 , n3251 );
not ( n11797 , n10472 );
nand ( n11798 , n11797 , n9089 );
nand ( n11799 , n7809 , n11798 );
and ( n11800 , n11799 , n7918 , n570 );
nor ( n11801 , n11796 , n11800 );
nor ( n11802 , n20 , n3493 , n6834 );
nor ( n11803 , n1387 , n11392 );
nand ( n11804 , n11803 , n10318 , n10683 , n10686 );
and ( n11805 , n7809 , n11804 );
or ( n11806 , n11510 , n11805 );
nand ( n11807 , n43 , n10687 );
or ( n11808 , n21 , n11807 );
nand ( n11809 , n11806 , n11808 , n11413 );
nand ( n11810 , n11802 , n11809 );
and ( n11811 , n11794 , n11801 , n11810 );
not ( n11812 , n20 );
not ( n11813 , n11738 );
nand ( n11814 , n7809 , n10654 );
not ( n11815 , n11814 );
or ( n11816 , n11813 , n11815 );
nand ( n11817 , n11816 , n11749 );
and ( n11818 , n11812 , n11817 );
nor ( n11819 , n571 , n11510 );
and ( n11820 , n11819 , n11799 );
nor ( n11821 , n628 , n11516 );
nor ( n11822 , n11820 , n11821 );
not ( n11823 , n11822 );
nor ( n11824 , n11818 , n11823 );
and ( n11825 , n11538 , n11673 );
nor ( n11826 , n11412 , n571 );
nand ( n11827 , n11826 , n10472 );
not ( n11828 , n11827 );
not ( n11829 , n16 );
nor ( n11830 , n7809 , n11829 , n630 );
nor ( n11831 , n11825 , n11828 , n11830 );
nand ( n11832 , n7809 , n10608 );
and ( n11833 , n11679 , n3146 , n11832 );
and ( n11834 , n2242 , n2446 );
nor ( n11835 , n11834 , n11537 );
nor ( n11836 , n11833 , n11835 );
and ( n11837 , n11538 , n2679 );
and ( n11838 , n11420 , n11814 );
not ( n11839 , n21 );
and ( n11840 , n43 , n10589 );
and ( n11841 , n11839 , n11840 );
nor ( n11842 , n11838 , n11841 );
and ( n11843 , n11413 , n11842 );
nor ( n11844 , n11843 , n6283 );
nor ( n11845 , n11837 , n11844 );
and ( n11846 , n11824 , n11831 , n11836 , n11845 );
and ( n11847 , n11766 , n11679 , n2515 );
not ( n11848 , n11805 );
and ( n11849 , n11848 , n11679 , n2243 );
nor ( n11850 , n11847 , n11849 );
not ( n11851 , n11777 );
not ( n11852 , n11851 );
and ( n11853 , n11852 , n11679 , n2679 );
and ( n11854 , n11420 , n11832 );
not ( n11855 , n21 );
not ( n11856 , n10198 );
nor ( n11857 , n7809 , n11856 );
and ( n11858 , n11855 , n11857 );
nor ( n11859 , n11854 , n11858 );
and ( n11860 , n11413 , n11859 );
not ( n11861 , n20 );
not ( n11862 , n3493 );
nand ( n11863 , n11861 , n11862 , n3299 );
nor ( n11864 , n11860 , n11863 );
nor ( n11865 , n11853 , n11864 );
nand ( n11866 , n11811 , n11846 , n11850 , n11865 );
or ( n11867 , n11782 , n11866 );
not ( n11868 , n18 );
nand ( n11869 , n11867 , n11868 );
not ( n11870 , n18 );
not ( n11871 , n11739 );
and ( n11872 , n11871 , n11394 );
and ( n11873 , n11712 , n11401 );
nor ( n11874 , n11872 , n11873 );
nand ( n11875 , n11874 , n11512 , n11518 );
not ( n11876 , n11714 );
not ( n11877 , n11408 );
or ( n11878 , n11876 , n11877 );
nand ( n11879 , n11878 , n11752 );
nor ( n11880 , n11875 , n11879 , n11431 , n11459 );
or ( n11881 , n11733 , n11546 );
or ( n11882 , n11725 , n11450 );
nand ( n11883 , n11881 , n11882 );
nand ( n11884 , n11526 , n11031 );
not ( n11885 , n11548 );
and ( n11886 , n11884 , n11885 );
nor ( n11887 , n11886 , n11428 , n6726 );
nor ( n11888 , n11883 , n11468 , n11887 );
and ( n11889 , n11735 , n11530 );
and ( n11890 , n11716 , n11443 );
nor ( n11891 , n11889 , n11890 );
not ( n11892 , n11526 );
not ( n11893 , n10793 );
or ( n11894 , n11892 , n11893 );
not ( n11895 , n11533 );
nand ( n11896 , n11894 , n11895 );
and ( n11897 , n11729 , n11896 );
or ( n11898 , n11412 , n11440 );
nand ( n11899 , n11898 , n11478 );
and ( n11900 , n11470 , n11899 );
nor ( n11901 , n11897 , n11900 );
nand ( n11902 , n11880 , n11888 , n11891 , n11901 );
and ( n11903 , n11870 , n11902 );
not ( n11904 , n11099 );
not ( n11905 , n10265 );
or ( n11906 , n11904 , n11905 );
nand ( n11907 , n11906 , n7809 );
and ( n11908 , n11738 , n11907 );
and ( n11909 , n11538 , n2816 );
nor ( n11910 , n11908 , n11909 , n11748 );
not ( n11911 , n10653 );
not ( n11912 , n10376 );
or ( n11913 , n11911 , n11912 );
nand ( n11914 , n11913 , n7809 );
and ( n11915 , n11420 , n11914 );
not ( n11916 , n10376 );
and ( n11917 , n11526 , n11916 );
nor ( n11918 , n11915 , n11917 );
and ( n11919 , n11413 , n11918 );
nor ( n11920 , n11919 , n3493 );
and ( n11921 , n11721 , n11920 );
or ( n11922 , n11537 , n11429 );
nand ( n11923 , n11922 , n11504 );
nor ( n11924 , n11921 , n11923 );
nand ( n11925 , n7809 , n11168 );
and ( n11926 , n11679 , n3299 , n11925 );
and ( n11927 , n11167 , n10320 );
nor ( n11928 , n11927 , n43 );
not ( n11929 , n11928 );
nand ( n11930 , n2816 , n11679 , n14 , n11929 );
not ( n11931 , n14 );
nand ( n11932 , n2816 , n11679 , n11931 , n11914 );
nand ( n11933 , n11930 , n11932 );
nor ( n11934 , n11926 , n11933 );
nand ( n11935 , n43 , n10200 );
or ( n11936 , n21 , n11935 );
not ( n11937 , n11925 );
or ( n11938 , n11510 , n11937 );
nand ( n11939 , n11936 , n11938 , n11413 );
not ( n11940 , n3516 );
and ( n11941 , n11939 , n11940 , n3299 );
and ( n11942 , n11420 , n11907 );
not ( n11943 , n21 );
nor ( n11944 , n7809 , n10265 );
and ( n11945 , n11943 , n11944 );
nor ( n11946 , n11942 , n11945 , n11477 );
or ( n11947 , n795 , n11946 );
or ( n11948 , n11510 , n11928 );
nand ( n11949 , n43 , n10406 );
or ( n11950 , n21 , n11949 );
nand ( n11951 , n11948 , n11950 , n11413 );
not ( n11952 , n3493 );
nand ( n11953 , n11951 , n11952 , n6835 );
nand ( n11954 , n11947 , n11953 );
nor ( n11955 , n11941 , n11954 );
nand ( n11956 , n11910 , n11924 , n11934 , n11955 );
and ( n11957 , n309 , n11956 );
not ( n11958 , n11819 );
not ( n11959 , n11670 );
or ( n11960 , n11958 , n11959 );
not ( n11961 , n9422 );
and ( n11962 , n11826 , n11961 );
nor ( n11963 , n11962 , n11821 );
nand ( n11964 , n11960 , n11963 );
and ( n11965 , n18 , n11964 );
nor ( n11966 , n11903 , n11957 , n11965 );
nand ( n11967 , n11710 , n11756 , n11869 , n11966 );
nand ( n11968 , n11967 , n4158 , n9012 );
nand ( n11969 , n1971 , n4241 , n4249 , n11967 );
and ( n11970 , n11664 , n11668 , n11968 , n11969 );
not ( n11971 , n21 );
and ( n11972 , n43 , n10498 );
and ( n11973 , n11971 , n11972 );
nor ( n11974 , n11973 , n11791 );
or ( n11975 , n11784 , n11974 );
and ( n11976 , n11538 , n10506 );
not ( n11977 , n3493 );
not ( n11978 , n11526 );
not ( n11979 , n10506 );
or ( n11980 , n11978 , n11979 );
nand ( n11981 , n11980 , n11768 );
nand ( n11982 , n11977 , n11981 );
not ( n11983 , n11982 );
or ( n11984 , n11398 , n11765 );
nand ( n11985 , n11984 , n11497 );
nor ( n11986 , n11976 , n11983 , n11985 );
or ( n11987 , n3128 , n11986 );
and ( n11988 , n11538 , n10762 );
and ( n11989 , n11397 , n11777 );
nor ( n11990 , n11989 , n11498 );
not ( n11991 , n11990 );
nand ( n11992 , n11526 , n10762 );
and ( n11993 , n11992 , n11779 );
nor ( n11994 , n11993 , n3493 );
nor ( n11995 , n11988 , n11991 , n11994 );
or ( n11996 , n2678 , n11995 );
nand ( n11997 , n11975 , n11987 , n11996 );
not ( n11998 , n11997 );
nor ( n11999 , n11482 , n2467 );
and ( n12000 , n11999 , n11972 );
nor ( n12001 , n20 , n11482 );
nand ( n12002 , n12001 , n6835 );
or ( n12003 , n12002 , n11807 );
nand ( n12004 , n12003 , n11810 );
nor ( n12005 , n11805 , n2242 , n11398 );
nor ( n12006 , n12000 , n12004 , n12005 );
and ( n12007 , n43 , n3345 , n10467 );
nor ( n12008 , n12007 , n11844 );
nand ( n12009 , n3146 , n11397 );
not ( n12010 , n12009 );
and ( n12011 , n12010 , n11832 );
nor ( n12012 , n20 , n11390 );
and ( n12013 , n12012 , n11814 );
nor ( n12014 , n12011 , n12013 );
not ( n12015 , n17 );
or ( n12016 , n12015 , n2242 );
nand ( n12017 , n12016 , n3346 );
and ( n12018 , n11492 , n12017 );
and ( n12019 , n11498 , n2468 );
not ( n12020 , n20 );
and ( n12021 , n12020 , n11505 );
nor ( n12022 , n12018 , n12019 , n12021 );
and ( n12023 , n12008 , n12014 , n11827 , n12022 );
nand ( n12024 , n3278 , n11840 );
not ( n12025 , n12024 );
not ( n12026 , n12001 );
nor ( n12027 , n7809 , n11429 );
not ( n12028 , n12027 );
or ( n12029 , n11856 , n12026 , n12028 );
nand ( n12030 , n3251 , n11397 );
or ( n12031 , n12030 , n11789 );
nand ( n12032 , n12029 , n12031 );
nand ( n12033 , n11389 , n570 );
not ( n12034 , n11799 );
or ( n12035 , n12033 , n12034 );
nand ( n12036 , n12035 , n11822 );
nor ( n12037 , n12025 , n12032 , n12036 , n11864 );
nand ( n12038 , n11998 , n12006 , n12023 , n12037 );
and ( n12039 , n11386 , n12038 );
and ( n12040 , n11999 , n11698 );
and ( n12041 , n12012 , n11907 );
nor ( n12042 , n12040 , n12041 );
not ( n12043 , n12042 );
or ( n12044 , n12009 , n11937 );
not ( n12045 , n11784 );
or ( n12046 , n11412 , n9471 );
nand ( n12047 , n12046 , n11701 );
and ( n12048 , n12045 , n12047 );
and ( n12049 , n11802 , n11951 );
nor ( n12050 , n12048 , n12049 );
nand ( n12051 , n12044 , n12050 );
not ( n12052 , n9545 );
and ( n12053 , n11538 , n12052 );
nand ( n12054 , n11526 , n9544 );
not ( n12055 , n11692 );
and ( n12056 , n12054 , n12055 );
nor ( n12057 , n12056 , n2781 );
not ( n12058 , n11397 );
not ( n12059 , n11689 );
or ( n12060 , n12058 , n12059 );
nand ( n12061 , n12060 , n11497 );
nor ( n12062 , n12053 , n12057 , n12061 );
or ( n12063 , n3128 , n12062 );
not ( n12064 , n11916 );
not ( n12065 , n12064 );
and ( n12066 , n11538 , n12065 );
and ( n12067 , n11397 , n11914 );
nor ( n12068 , n12067 , n11498 );
not ( n12069 , n11920 );
nand ( n12070 , n12068 , n12069 );
nor ( n12071 , n12066 , n12070 );
or ( n12072 , n2678 , n12071 );
and ( n12073 , n10200 , n12001 , n12027 );
not ( n12074 , n11863 );
and ( n12075 , n12074 , n11939 );
nor ( n12076 , n12073 , n12075 );
nand ( n12077 , n12063 , n12072 , n12076 );
or ( n12078 , n12002 , n11949 );
nand ( n12079 , n3278 , n11944 );
nand ( n12080 , n12078 , n12079 );
nor ( n12081 , n12043 , n12051 , n12077 , n12080 );
not ( n12082 , n12033 );
not ( n12083 , n11670 );
not ( n12084 , n12083 );
and ( n12085 , n12082 , n12084 );
not ( n12086 , n11964 );
nand ( n12087 , n12086 , n12022 );
nor ( n12088 , n12085 , n12087 );
and ( n12089 , n11929 , n2243 , n11397 );
and ( n12090 , n11830 , n11961 );
nor ( n12091 , n12089 , n12090 );
not ( n12092 , n6283 );
not ( n12093 , n11946 );
and ( n12094 , n12092 , n12093 );
not ( n12095 , n11681 );
nor ( n12096 , n12030 , n12095 );
nor ( n12097 , n12094 , n12096 );
nand ( n12098 , n12081 , n12088 , n12091 , n12097 );
and ( n12099 , n11560 , n12098 );
nor ( n12100 , n12039 , n12099 );
not ( n12101 , n8622 );
not ( n12102 , n12101 );
not ( n12103 , n12102 );
not ( n12104 , n12103 );
not ( n12105 , n12104 );
not ( n12106 , n12105 );
not ( n12107 , n12106 );
not ( n12108 , n12107 );
and ( n12109 , n12108 , n10958 );
nor ( n12110 , n12109 , n11409 );
not ( n12111 , n12110 );
nor ( n12112 , n31 , n2898 );
or ( n12113 , n7809 , n12112 );
nand ( n12114 , n12111 , n12113 );
and ( n12115 , n1419 , n12114 );
and ( n12116 , n1371 , n1409 );
nand ( n12117 , n43 , n5103 );
nor ( n12118 , n12116 , n12117 );
nor ( n12119 , n12115 , n12118 );
nand ( n12120 , n10465 , n11602 );
not ( n12121 , n10466 );
not ( n12122 , n10464 );
nor ( n12123 , n12120 , n12121 , n12122 );
or ( n12124 , n12123 , n12034 );
nand ( n12125 , n12124 , n12113 );
and ( n12126 , n12125 , n1370 , n1374 );
not ( n12127 , n8631 );
and ( n12128 , n12127 , n6762 );
nor ( n12129 , n12128 , n12117 );
nor ( n12130 , n12126 , n12129 );
not ( n12131 , n12120 );
and ( n12132 , n12131 , n9605 , n10838 , n10841 );
not ( n12133 , n11443 );
or ( n12134 , n12132 , n12133 );
nand ( n12135 , n12134 , n12113 );
and ( n12136 , n12135 , n1406 , n764 );
not ( n12137 , n12108 );
or ( n12138 , n12137 , n11050 );
nand ( n12139 , n12138 , n11545 );
nand ( n12140 , n12113 , n12139 );
and ( n12141 , n1909 , n12140 );
nor ( n12142 , n12136 , n12141 );
not ( n12143 , n3451 );
nand ( n12144 , n12131 , n10318 , n10683 , n10686 );
and ( n12145 , n12144 , n11848 );
not ( n12146 , n12113 );
nor ( n12147 , n12145 , n12146 );
not ( n12148 , n12147 );
and ( n12149 , n12143 , n12148 );
nand ( n12150 , n12131 , n9911 , n10890 , n10892 );
and ( n12151 , n12150 , n11449 );
nor ( n12152 , n12151 , n12146 );
nor ( n12153 , n1913 , n12152 );
nor ( n12154 , n12149 , n12153 );
nand ( n12155 , n12119 , n12130 , n12142 , n12154 );
and ( n12156 , n12103 , n11832 );
nor ( n12157 , n12156 , n12146 , n11857 );
or ( n12158 , n1612 , n12157 );
not ( n12159 , n10589 );
nand ( n12160 , n12159 , n12104 );
and ( n12161 , n12160 , n11814 );
nor ( n12162 , n12161 , n12146 );
or ( n12163 , n1143 , n12162 );
or ( n12164 , n12105 , n10923 );
nand ( n12165 , n12164 , n11530 );
nand ( n12166 , n12113 , n12165 );
and ( n12167 , n12166 , n1406 , n583 );
and ( n12168 , n12131 , n9469 , n10495 , n10497 );
or ( n12169 , n12168 , n11789 );
nand ( n12170 , n12169 , n12113 );
and ( n12171 , n1787 , n12170 );
nor ( n12172 , n12167 , n12171 );
nand ( n12173 , n12158 , n12163 , n12172 );
nand ( n12174 , n12108 , n10987 );
and ( n12175 , n12174 , n11394 );
nor ( n12176 , n12175 , n12146 );
or ( n12177 , n1947 , n12176 );
not ( n12178 , n12137 );
nand ( n12179 , n12178 , n10851 );
and ( n12180 , n12179 , n11401 );
nor ( n12181 , n12180 , n12146 );
or ( n12182 , n1941 , n12181 );
not ( n12183 , n10505 );
or ( n12184 , n12103 , n12183 );
nand ( n12185 , n12184 , n11766 );
nand ( n12186 , n12113 , n12185 );
and ( n12187 , n1432 , n12186 );
nand ( n12188 , n12131 , n10336 , n10751 , n10754 );
and ( n12189 , n12188 , n11777 );
nor ( n12190 , n12189 , n12146 );
not ( n12191 , n12190 );
and ( n12192 , n1223 , n12191 );
nor ( n12193 , n12187 , n12192 );
nand ( n12194 , n12177 , n12182 , n12193 );
nor ( n12195 , n12155 , n12173 , n12194 );
or ( n12196 , n3748 , n12195 );
not ( n12197 , n7809 );
not ( n12198 , n11604 );
and ( n12199 , n12197 , n12198 );
nor ( n12200 , n12199 , n12146 );
nor ( n12201 , n3748 , n12200 );
and ( n12202 , n12201 , n3425 , n724 );
not ( n12203 , n3748 );
and ( n12204 , n43 , n11589 );
or ( n12205 , n12146 , n12204 );
and ( n12206 , n12203 , n2003 , n12205 );
nor ( n12207 , n12202 , n12206 );
not ( n12208 , n12207 );
nor ( n12209 , n3747 , n1989 );
nor ( n12210 , n11603 , n9307 );
or ( n12211 , n7809 , n12210 );
nand ( n12212 , n12211 , n12113 );
and ( n12213 , n12209 , n12212 );
nor ( n12214 , n7809 , n12102 );
nor ( n12215 , n11944 , n12146 , n12214 );
or ( n12216 , n3928 , n6283 , n12215 );
nor ( n12217 , n11629 , n12146 , n12214 );
or ( n12218 , n3747 , n2022 , n12217 );
nand ( n12219 , n12216 , n12218 );
not ( n12220 , n96 );
not ( n12221 , n12105 );
and ( n12222 , n12221 , n9975 );
nor ( n12223 , n12222 , n11659 );
nor ( n12224 , n12146 , n12223 );
nor ( n12225 , n12220 , n3747 , n12224 , n1599 );
nor ( n12226 , n12213 , n12219 , n12225 );
nor ( n12227 , n12117 , n3747 );
and ( n12228 , n9038 , n12227 );
and ( n12229 , n43 , n3748 );
nor ( n12230 , n12228 , n12229 );
or ( n12231 , n9591 , n2863 );
nand ( n12232 , n12231 , n12227 );
not ( n12233 , n1583 );
or ( n12234 , n2009 , n12233 );
nand ( n12235 , n12234 , n12227 );
nand ( n12236 , n12226 , n12230 , n12232 , n12235 );
nand ( n12237 , n12106 , n9607 );
and ( n12238 , n12237 , n11562 );
nor ( n12239 , n12238 , n12146 );
or ( n12240 , n12239 , n632 , n9108 );
not ( n12241 , n3748 );
nor ( n12242 , n8621 , n11961 );
or ( n12243 , n12242 , n12083 );
nand ( n12244 , n12243 , n12113 );
nand ( n12245 , n309 , n12241 , n1374 , n12244 );
nand ( n12246 , n12240 , n12245 );
not ( n12247 , n12103 );
nand ( n12248 , n12247 , n10407 );
and ( n12249 , n12248 , n11929 );
nor ( n12250 , n12249 , n12146 );
or ( n12251 , n12250 , n3928 , n6286 );
nand ( n12252 , n12102 , n9708 );
not ( n12253 , n11566 );
and ( n12254 , n12252 , n12253 );
nor ( n12255 , n12254 , n12146 );
or ( n12256 , n12255 , n521 , n9108 );
nand ( n12257 , n12251 , n12256 );
nor ( n12258 , n12208 , n12236 , n12246 , n12257 );
nand ( n12259 , n12196 , n12258 );
nand ( n12260 , n3787 , n2617 );
nand ( n12261 , n12104 , n12064 );
and ( n12262 , n12261 , n11914 );
nor ( n12263 , n12262 , n12146 );
or ( n12264 , n12260 , n12263 );
not ( n12265 , n3748 );
not ( n12266 , n1581 );
or ( n12267 , n8621 , n9470 );
nand ( n12268 , n12267 , n11681 );
nand ( n12269 , n12113 , n12268 );
nand ( n12270 , n590 , n12265 , n12266 , n12269 );
nand ( n12271 , n12264 , n12270 );
and ( n12272 , n12107 , n11925 );
nand ( n12273 , n12113 , n11935 );
nor ( n12274 , n12272 , n12273 );
or ( n12275 , n12274 , n3928 , n3264 );
nand ( n12276 , n309 , n583 );
or ( n12277 , n11603 , n9542 );
nand ( n12278 , n12277 , n11689 );
nand ( n12279 , n12113 , n12278 );
not ( n12280 , n12279 );
or ( n12281 , n12276 , n3748 , n12280 );
nand ( n12282 , n12275 , n12281 );
or ( n12283 , n12259 , n12271 , n12282 );
nand ( n12284 , n12283 , n4258 );
not ( n12285 , n3748 );
nor ( n12286 , n18 , n1 , n12285 );
and ( n12287 , n2418 , n11814 );
not ( n12288 , n20 );
not ( n12289 , n3493 );
and ( n12290 , n12289 , n2937 );
nor ( n12291 , n12290 , n7809 );
and ( n12292 , n12288 , n12291 );
nor ( n12293 , n12287 , n12292 );
and ( n12294 , n3281 , n11832 );
and ( n12295 , n2463 , n11799 );
nor ( n12296 , n12294 , n12295 );
not ( n12297 , n3417 );
not ( n12298 , n11805 );
and ( n12299 , n12297 , n12298 );
and ( n12300 , n3413 , n11795 );
nor ( n12301 , n12299 , n12300 );
and ( n12302 , n3350 , n11766 );
and ( n12303 , n3025 , n11852 );
nor ( n12304 , n12302 , n12303 );
nand ( n12305 , n12293 , n12296 , n12301 , n12304 );
and ( n12306 , n12286 , n12305 );
and ( n12307 , n2544 , n11408 );
and ( n12308 , n20 , n12291 );
nor ( n12309 , n12307 , n12308 );
and ( n12310 , n11443 , n908 , n2736 );
not ( n12311 , n11401 );
nor ( n12312 , n2551 , n12311 );
nor ( n12313 , n12310 , n12312 );
and ( n12314 , n2304 , n11545 );
and ( n12315 , n3221 , n11394 );
nor ( n12316 , n12314 , n12315 );
and ( n12317 , n3399 , n11530 );
and ( n12318 , n2559 , n11449 );
nor ( n12319 , n12317 , n12318 );
nand ( n12320 , n12309 , n12313 , n12316 , n12319 );
and ( n12321 , n12286 , n12320 );
nor ( n12322 , n12306 , n12321 );
not ( n12323 , n12322 );
not ( n12324 , n11907 );
nor ( n12325 , n1 , n20 );
nand ( n12326 , n18 , n12325 );
nand ( n12327 , n3748 , n2802 );
or ( n12328 , n12324 , n12326 , n12327 );
not ( n12329 , n18 );
nor ( n12330 , n12329 , n1 );
nand ( n12331 , n12330 , n3748 , n2463 , n11670 );
nand ( n12332 , n12328 , n12331 );
not ( n12333 , n9496 );
nor ( n12334 , n12333 , n1 );
nand ( n12335 , n12334 , n522 );
not ( n12336 , n3748 );
or ( n12337 , n12335 , n12336 , n11707 );
nand ( n12338 , n2506 , n1582 );
or ( n12339 , n11625 , n12338 , n12327 );
nand ( n12340 , n12337 , n12339 );
not ( n12341 , n11914 );
nand ( n12342 , n3748 , n2800 );
or ( n12343 , n12341 , n12326 , n12342 );
nand ( n12344 , n3748 , n11644 );
or ( n12345 , n12344 , n12338 , n2791 );
nand ( n12346 , n12343 , n12345 );
nor ( n12347 , n12323 , n12332 , n12340 , n12346 );
not ( n12348 , n12330 );
not ( n12349 , n2195 );
or ( n12350 , n12348 , n12349 );
or ( n12351 , n1 , n1575 );
nand ( n12352 , n12350 , n12351 );
and ( n12353 , n12352 , n3748 , n12291 );
not ( n12354 , n19 );
and ( n12355 , n12354 , n12291 );
and ( n12356 , n12355 , n12330 , n3748 );
nor ( n12357 , n12353 , n12356 );
nand ( n12358 , n11288 , n2544 , n2506 , n11578 );
nand ( n12359 , n12330 , n3748 , n3413 , n11681 );
nand ( n12360 , n12347 , n12357 , n12358 , n12359 );
nand ( n12361 , n12330 , n2489 , n3748 , n11562 );
not ( n12362 , n12326 );
not ( n12363 , n3748 );
nor ( n12364 , n12363 , n2789 );
nand ( n12365 , n12362 , n11929 , n12364 );
not ( n12366 , n12338 );
nand ( n12367 , n12366 , n11635 , n12364 );
nand ( n12368 , n12325 , n11288 , n2538 , n11925 );
nand ( n12369 , n12361 , n12365 , n12367 , n12368 );
not ( n12370 , n3748 );
nand ( n12371 , n2506 , n12370 );
nand ( n12372 , n43 , n2303 );
and ( n12373 , n12110 , n12372 , n1921 );
not ( n12374 , n448 );
nor ( n12375 , n7809 , n12374 );
and ( n12376 , n16 , n12375 );
nor ( n12377 , n2744 , n12113 );
and ( n12378 , n7039 , n12377 );
nor ( n12379 , n12376 , n12378 );
and ( n12380 , n6674 , n12377 );
not ( n12381 , n14 );
not ( n12382 , n16 );
nand ( n12383 , n12381 , n12382 );
nor ( n12384 , n2303 , n12383 );
and ( n12385 , n12384 , n12146 );
not ( n12386 , n16 );
and ( n12387 , n12386 , n12375 );
nor ( n12388 , n12380 , n12385 , n12387 );
and ( n12389 , n12379 , n12388 );
nor ( n12390 , n12389 , n1315 );
nor ( n12391 , n12373 , n12390 );
not ( n12392 , n18 );
and ( n12393 , n12392 , n7695 , n12114 );
nand ( n12394 , n2303 , n1314 );
nor ( n12395 , n12176 , n521 , n12394 );
nor ( n12396 , n12393 , n12395 );
not ( n12397 , n18 );
nand ( n12398 , n12397 , n7809 , n2409 , n11408 );
and ( n12399 , n43 , n2744 );
nor ( n12400 , n12399 , n7038 );
nand ( n12401 , n1314 , n12400 , n11423 );
and ( n12402 , n12391 , n12396 , n12398 , n12401 );
not ( n12403 , n12102 );
not ( n12404 , n12372 );
nor ( n12405 , n12404 , n12383 );
and ( n12406 , n12403 , n12405 );
nor ( n12407 , n43 , n2498 );
nor ( n12408 , n12406 , n12407 );
not ( n12409 , n12408 );
and ( n12410 , n12409 , n11394 );
and ( n12411 , n12405 , n11455 );
nor ( n12412 , n12410 , n12411 );
or ( n12413 , n1315 , n12412 );
not ( n12414 , n12399 );
not ( n12415 , n8617 );
and ( n12416 , n12414 , n12415 );
nor ( n12417 , n43 , n2744 );
nor ( n12418 , n12416 , n12417 );
nor ( n12419 , n7038 , n12418 );
and ( n12420 , n11401 , n1314 , n12419 );
nor ( n12421 , n2303 , n12113 );
or ( n12422 , n12375 , n12421 );
and ( n12423 , n1921 , n12422 );
nor ( n12424 , n12420 , n12423 );
nand ( n12425 , n12413 , n12424 );
nand ( n12426 , n1317 , n11545 );
or ( n12427 , n12426 , n2303 , n43 );
not ( n12428 , n11183 );
or ( n12429 , n12399 , n12428 , n11461 );
nand ( n12430 , n12427 , n12429 );
nor ( n12431 , n11450 , n12428 , n12418 );
nand ( n12432 , n8026 , n7039 );
not ( n12433 , n12432 );
and ( n12434 , n12433 , n12135 );
and ( n12435 , n12419 , n11443 );
and ( n12436 , n12400 , n11473 );
nor ( n12437 , n12434 , n12435 , n12436 );
nor ( n12438 , n42 , n521 );
and ( n12439 , n12438 , n12166 );
nor ( n12440 , n12387 , n12378 );
not ( n12441 , n12440 );
nor ( n12442 , n12439 , n12441 );
and ( n12443 , n12384 , n11541 );
and ( n12444 , n12407 , n11530 );
nor ( n12445 , n12443 , n12444 );
and ( n12446 , n12437 , n12442 , n12445 );
nor ( n12447 , n12446 , n1415 );
nor ( n12448 , n12425 , n12430 , n12431 , n12447 );
not ( n12449 , n12394 );
and ( n12450 , n12140 , n724 , n12449 );
nor ( n12451 , n12181 , n1315 , n12432 );
nor ( n12452 , n12450 , n12451 );
nor ( n12453 , n12152 , n2937 , n12428 );
not ( n12454 , n18 );
not ( n12455 , n12454 );
and ( n12456 , n8044 , n12372 , n12101 );
and ( n12457 , n7809 , n2802 );
nor ( n12458 , n12456 , n12457 );
nor ( n12459 , n20 , n12458 );
and ( n12460 , n12459 , n11814 );
not ( n12461 , n12024 );
and ( n12462 , n12372 , n12461 );
nor ( n12463 , n12460 , n12462 );
or ( n12464 , n6676 , n11157 );
nand ( n12465 , n12464 , n12377 );
and ( n12466 , n12375 , n3256 );
and ( n12467 , n453 , n12376 );
and ( n12468 , n3278 , n12421 );
nor ( n12469 , n12466 , n12467 , n12468 );
nand ( n12470 , n12463 , n12465 , n12469 );
not ( n12471 , n11832 );
or ( n12472 , n12418 , n11243 , n12471 );
nand ( n12473 , n8026 , n11157 );
or ( n12474 , n12473 , n12157 );
nand ( n12475 , n12472 , n12474 );
nand ( n12476 , n2303 , n2255 );
or ( n12477 , n12476 , n12190 );
nand ( n12478 , n2303 , n2417 );
or ( n12479 , n12478 , n12162 );
nand ( n12480 , n12477 , n12479 );
nor ( n12481 , n12470 , n12475 , n12480 );
not ( n12482 , n12418 );
and ( n12483 , n11848 , n6676 , n12482 );
not ( n12484 , n19 );
nand ( n12485 , n12484 , n15 , n2998 );
or ( n12486 , n12147 , n6675 , n12485 );
not ( n12487 , n14 );
nand ( n12488 , n12487 , n2816 , n2461 );
or ( n12489 , n11482 , n11774 );
nand ( n12490 , n12489 , n11990 );
nor ( n12491 , n12490 , n11994 );
or ( n12492 , n12488 , n12491 );
nand ( n12493 , n12486 , n12492 );
nor ( n12494 , n12483 , n12493 );
not ( n12495 , n12399 );
nand ( n12496 , n12495 , n6676 );
not ( n12497 , n12496 );
not ( n12498 , n11807 );
and ( n12499 , n12497 , n12498 );
nor ( n12500 , n12399 , n11243 );
and ( n12501 , n12500 , n11857 );
nor ( n12502 , n12499 , n12501 );
not ( n12503 , n20 );
nor ( n12504 , n43 , n3349 );
and ( n12505 , n12504 , n11766 );
nor ( n12506 , n42 , n1375 );
not ( n12507 , n12506 );
not ( n12508 , n12125 );
or ( n12509 , n12507 , n12508 );
and ( n12510 , n1373 , n12372 , n8620 );
and ( n12511 , n7809 , n42 , n1374 );
nor ( n12512 , n12510 , n12511 );
not ( n12513 , n12512 );
and ( n12514 , n12513 , n11799 );
nor ( n12515 , n7809 , n1372 , n12404 );
and ( n12516 , n12515 , n10472 );
nor ( n12517 , n12514 , n12516 );
nand ( n12518 , n12509 , n12517 );
nor ( n12519 , n11076 , n12418 );
not ( n12520 , n12519 );
or ( n12521 , n12520 , n11789 );
and ( n12522 , n1373 , n12422 );
and ( n12523 , n11075 , n12377 );
and ( n12524 , n19 , n12387 );
nor ( n12525 , n12522 , n12523 , n12524 );
nand ( n12526 , n12521 , n12525 );
nor ( n12527 , n12505 , n12518 , n12526 );
nor ( n12528 , n42 , n1880 );
and ( n12529 , n12528 , n12186 );
nor ( n12530 , n12399 , n11076 );
and ( n12531 , n12530 , n11972 );
nor ( n12532 , n12529 , n12531 );
not ( n12533 , n19 );
nor ( n12534 , n12533 , n2937 );
and ( n12535 , n12170 , n7039 , n12534 );
and ( n12536 , n11483 , n11760 );
nor ( n12537 , n12536 , n11985 );
and ( n12538 , n12537 , n11982 );
nand ( n12539 , n19 , n12384 );
nor ( n12540 , n12538 , n12539 );
nor ( n12541 , n12535 , n12540 );
nand ( n12542 , n12527 , n12532 , n12541 );
and ( n12543 , n12503 , n12542 );
nand ( n12544 , n7809 , n453 , n3426 );
nor ( n12545 , n12544 , n11851 );
nor ( n12546 , n12543 , n12545 );
nand ( n12547 , n12481 , n12494 , n12502 , n12546 );
not ( n12548 , n12547 );
or ( n12549 , n12455 , n12548 );
not ( n12550 , n16 );
nor ( n12551 , n12550 , n14 );
nand ( n12552 , n12551 , n42 , n1314 , n11554 );
nand ( n12553 , n12549 , n12552 );
nor ( n12554 , n12453 , n12553 );
and ( n12555 , n12402 , n12448 , n12452 , n12554 );
or ( n12556 , n12371 , n12555 );
not ( n12557 , n3748 );
nor ( n12558 , n12557 , n11566 );
and ( n12559 , n12558 , n12334 , n909 );
nor ( n12560 , n43 , n11600 );
and ( n12561 , n12560 , n3425 , n3426 );
nor ( n12562 , n11659 , n11091 , n12418 );
nor ( n12563 , n12561 , n12562 );
or ( n12564 , n1599 , n12388 );
and ( n12565 , n18 , n7695 , n12212 );
and ( n12566 , n1975 , n12422 );
nor ( n12567 , n12565 , n12566 );
nand ( n12568 , n12564 , n12567 );
or ( n12569 , n11625 , n1599 , n12408 );
not ( n12570 , n12210 );
and ( n12571 , n12570 , n12372 , n1975 );
and ( n12572 , n7809 , n18 , n2409 );
nor ( n12573 , n12571 , n12572 );
or ( n12574 , n11579 , n12573 );
nand ( n12575 , n12569 , n12574 );
nor ( n12576 , n7038 , n1599 );
and ( n12577 , n11644 , n12417 , n12576 );
nor ( n12578 , n12399 , n1599 );
and ( n12579 , n7039 , n12578 , n12204 );
nor ( n12580 , n12577 , n12579 );
not ( n12581 , n12580 );
nor ( n12582 , n12568 , n12575 , n12581 );
and ( n12583 , n8026 , n12576 , n12205 );
and ( n12584 , n12405 , n3425 , n11629 );
nor ( n12585 , n12583 , n12584 );
nor ( n12586 , n42 , n12200 );
and ( n12587 , n12586 , n3425 , n724 );
and ( n12588 , n6674 , n12578 , n11638 );
nor ( n12589 , n12587 , n12588 );
nand ( n12590 , n12563 , n12582 , n12585 , n12589 );
or ( n12591 , n12224 , n2937 , n11091 );
not ( n12592 , n12438 );
or ( n12593 , n12592 , n1599 , n12217 );
nand ( n12594 , n12591 , n12593 );
not ( n12595 , n11611 );
nand ( n12596 , n12595 , n42 , n3425 );
not ( n12597 , n16 );
or ( n12598 , n12596 , n12597 , n14 );
or ( n12599 , n1599 , n12379 );
nand ( n12600 , n12598 , n12599 );
nor ( n12601 , n12590 , n12594 , n12600 );
not ( n12602 , n12400 );
not ( n12603 , n11616 );
or ( n12604 , n12602 , n12603 );
and ( n12605 , n12419 , n11562 );
and ( n12606 , n12407 , n12253 );
nor ( n12607 , n12605 , n12606 );
nand ( n12608 , n12604 , n12607 );
or ( n12609 , n12432 , n12239 );
not ( n12610 , n11574 );
and ( n12611 , n12384 , n12610 );
not ( n12612 , n12255 );
and ( n12613 , n12438 , n12612 );
nor ( n12614 , n12611 , n12613 );
nand ( n12615 , n12609 , n12614 , n12440 );
or ( n12616 , n12608 , n12615 );
nand ( n12617 , n12616 , n3242 );
and ( n12618 , n12459 , n11907 );
not ( n12619 , n12469 );
nor ( n12620 , n12618 , n12619 );
nand ( n12621 , n12482 , n11157 , n11925 );
nand ( n12622 , n12620 , n12465 , n12621 );
or ( n12623 , n12478 , n12215 );
or ( n12624 , n2303 , n12079 );
nand ( n12625 , n12623 , n12624 );
or ( n12626 , n12250 , n6675 , n12485 );
or ( n12627 , n12544 , n12341 );
nand ( n12628 , n12626 , n12627 );
nor ( n12629 , n12622 , n12625 , n12628 );
and ( n12630 , n11929 , n6676 , n12482 );
and ( n12631 , n12515 , n11961 );
and ( n12632 , n12506 , n12244 );
or ( n12633 , n12512 , n12083 );
nand ( n12634 , n12504 , n11689 );
nand ( n12635 , n12633 , n12634 , n12525 );
nor ( n12636 , n12631 , n12632 , n12635 );
and ( n12637 , n12528 , n12279 );
and ( n12638 , n12519 , n11681 );
and ( n12639 , n12530 , n11698 );
nor ( n12640 , n12637 , n12638 , n12639 );
not ( n12641 , n12539 );
not ( n12642 , n11483 );
not ( n12643 , n11685 );
or ( n12644 , n12642 , n12643 );
not ( n12645 , n12061 );
nand ( n12646 , n12644 , n12645 );
nor ( n12647 , n12646 , n12057 );
not ( n12648 , n12647 );
and ( n12649 , n12641 , n12648 );
and ( n12650 , n12269 , n7039 , n12534 );
nor ( n12651 , n12649 , n12650 );
and ( n12652 , n12636 , n12640 , n12651 );
or ( n12653 , n20 , n12652 );
or ( n12654 , n12476 , n12263 );
nand ( n12655 , n12653 , n12654 );
nor ( n12656 , n12630 , n12655 );
not ( n12657 , n12496 );
not ( n12658 , n11949 );
and ( n12659 , n12657 , n12658 );
not ( n12660 , n12500 );
nor ( n12661 , n12660 , n11935 );
nor ( n12662 , n12659 , n12661 );
not ( n12663 , n12473 );
not ( n12664 , n12274 );
and ( n12665 , n12663 , n12664 );
nand ( n12666 , n43 , n11483 , n12065 );
and ( n12667 , n12068 , n12666 , n12069 );
nor ( n12668 , n12667 , n12488 );
nor ( n12669 , n12665 , n12668 );
nand ( n12670 , n12629 , n12656 , n12662 , n12669 );
nand ( n12671 , n18 , n12670 );
and ( n12672 , n12601 , n12617 , n12671 );
nor ( n12673 , n12672 , n12371 );
nor ( n12674 , n12559 , n12673 );
or ( n12675 , n11600 , n12338 , n12342 );
nand ( n12676 , n12556 , n12674 , n12675 );
or ( n12677 , n12360 , n12369 , n12676 );
nor ( n12678 , n4261 , n4240 );
nand ( n12679 , n12677 , n12678 );
nand ( n12680 , n11970 , n12100 , n12284 , n12679 );
or ( n12681 , n9014 , n4234 );
not ( n12682 , n7 );
nor ( n12683 , n12682 , n4234 );
and ( n12684 , n8 , n31 );
nand ( n12685 , n10 , n12684 );
not ( n12686 , n12685 );
and ( n12687 , n12683 , n12686 );
and ( n12688 , n7 , n12684 );
nor ( n12689 , n4236 , n7 );
nor ( n12690 , n12688 , n9 , n12689 );
nor ( n12691 , n12682 , n10 );
nor ( n12692 , n5820 , n10430 );
not ( n12693 , n12692 );
nand ( n12694 , n34 , n3815 );
nand ( n12695 , n12693 , n12694 );
and ( n12696 , n8 , n9 , n12691 , n12695 );
nor ( n12697 , n12687 , n12690 , n12696 );
and ( n12698 , n12 , n5315 , n8885 );
not ( n12699 , n8885 );
not ( n12700 , n40 );
not ( n12701 , n2 );
and ( n12702 , n13 , n12701 );
not ( n12703 , n12702 );
nor ( n12704 , n12699 , n12700 , n12 , n12703 );
nor ( n12705 , n12698 , n12704 );
not ( n12706 , n12705 );
not ( n12707 , n313 );
nand ( n12708 , n2309 , n12707 );
not ( n12709 , n12708 );
or ( n12710 , n8886 , n3838 , n12709 );
not ( n12711 , n23 );
nor ( n12712 , n12711 , n24 );
and ( n12713 , n12712 , n3762 );
and ( n12714 , n23 , n3812 );
not ( n12715 , n12714 );
not ( n12716 , n12715 );
not ( n12717 , n12716 );
nor ( n12718 , n12713 , n12717 );
not ( n12719 , n12718 );
nor ( n12720 , n4159 , n1852 );
nand ( n12721 , n12719 , n3753 , n12720 );
nand ( n12722 , n12710 , n12721 );
or ( n12723 , n2 , n13 );
nand ( n12724 , n12723 , n3523 );
or ( n12725 , n12724 , n5314 , n8886 );
not ( n12726 , n3753 );
nor ( n12727 , n12726 , n3761 );
nand ( n12728 , n4157 , n12727 );
nor ( n12729 , n2 , n12 );
not ( n12730 , n40 );
nand ( n12731 , n12730 , n5312 );
and ( n12732 , n13 , n12729 , n12731 );
not ( n12733 , n2 );
nand ( n12734 , n1845 , n12733 , n3837 );
not ( n12735 , n12734 );
not ( n12736 , n12735 );
not ( n12737 , n13 );
nand ( n12738 , n12737 , n12729 );
not ( n12739 , n12738 );
nand ( n12740 , n86 , n5312 );
nand ( n12741 , n12739 , n12740 );
nand ( n12742 , n12736 , n12741 );
nor ( n12743 , n12732 , n12742 );
or ( n12744 , n12728 , n12743 );
nand ( n12745 , n12725 , n12744 );
nand ( n12746 , n5897 , n12735 );
or ( n12747 , n3755 , n12746 );
not ( n12748 , n987 );
not ( n12749 , n24 );
not ( n12750 , n40 );
or ( n12751 , n12749 , n12750 );
nand ( n12752 , n12751 , n12714 );
not ( n12753 , n12752 );
or ( n12754 , n12748 , n12753 );
or ( n12755 , n445 , n12715 );
not ( n12756 , n24 );
nor ( n12757 , n12756 , n40 );
not ( n12758 , n12714 );
nor ( n12759 , n12757 , n12758 );
nand ( n12760 , n445 , n12759 );
nand ( n12761 , n12755 , n80 , n12760 );
nand ( n12762 , n12754 , n12761 );
not ( n12763 , n12762 );
and ( n12764 , n445 , n12715 );
not ( n12765 , n445 );
not ( n12766 , n12759 );
and ( n12767 , n12765 , n12766 );
nor ( n12768 , n12764 , n12767 );
not ( n12769 , n12768 );
nand ( n12770 , n3531 , n12769 );
not ( n12771 , n3520 );
nand ( n12772 , n1980 , n3524 );
not ( n12773 , n12772 );
not ( n12774 , n12773 );
or ( n12775 , n12771 , n12774 );
nand ( n12776 , n12715 , n7793 , n12734 );
nand ( n12777 , n12746 , n12776 );
nand ( n12778 , n12775 , n12777 );
nand ( n12779 , n12763 , n12770 , n12778 );
nand ( n12780 , n2888 , n4 , n12779 );
nand ( n12781 , n12747 , n12780 );
nor ( n12782 , n12706 , n12722 , n12745 , n12781 );
and ( n12783 , n8885 , n12742 );
nand ( n12784 , n3761 , n3753 );
not ( n12785 , n993 );
nor ( n12786 , n12785 , n3756 );
not ( n12787 , n12786 );
nor ( n12788 , n12718 , n12787 , n3755 );
nor ( n12789 , n12783 , t_0 , n12788 );
not ( n12790 , n12709 );
nand ( n12791 , n12790 , n12727 , n6440 );
not ( n12792 , n24 );
nand ( n12793 , n12792 , n39 );
not ( n12794 , n12715 );
nand ( n12795 , n12793 , n12794 );
nand ( n12796 , n5 , n994 , n4157 , n12795 );
nand ( n12797 , n5 , n3609 , n6440 , n12769 );
nand ( n12798 , n5 , n2298 );
nor ( n12799 , n2506 , n12798 );
not ( n12800 , n2 );
not ( n12801 , n3837 );
and ( n12802 , n12800 , n1845 , n12801 );
nand ( n12803 , n12 , n12795 , n12799 , n12802 );
nor ( n12804 , n2299 , n4015 );
nand ( n12805 , n12804 , n1852 , n2508 , n12769 );
nand ( n12806 , n12796 , n12797 , n12803 , n12805 );
nand ( n12807 , n5 , n4160 , n1852 , n12708 );
nor ( n12808 , n39 , n4174 );
nand ( n12809 , n12808 , n2508 , n1852 , n12708 );
not ( n12810 , n12798 );
not ( n12811 , n12712 );
not ( n12812 , n4013 );
or ( n12813 , n12811 , n12812 );
nand ( n12814 , n12813 , n12716 );
nand ( n12815 , n12810 , n2506 , n12814 , n12786 );
not ( n12816 , n12743 );
nand ( n12817 , n12816 , n2507 , n12808 );
nand ( n12818 , n12807 , n12809 , n12815 , n12817 );
nor ( n12819 , n12806 , n12818 );
not ( n12820 , n12799 );
not ( n12821 , n5899 );
or ( n12822 , n12820 , n12821 );
and ( n12823 , n1 , n5 );
nand ( n12824 , n39 , n2298 , n12823 );
nand ( n12825 , n12822 , n12824 );
and ( n12826 , n12735 , n12825 );
not ( n12827 , n12740 );
or ( n12828 , n12824 , n81 , n12827 );
nand ( n12829 , n12 , n12823 , n12795 );
not ( n12830 , n2 );
or ( n12831 , n12829 , n12830 , n3 );
nand ( n12832 , n12828 , n12831 );
not ( n12833 , n4187 );
not ( n12834 , n12779 );
or ( n12835 , n12833 , n12834 );
nand ( n12836 , n5 , n4158 , n3523 , n12795 );
nand ( n12837 , n12835 , n12836 );
nor ( n12838 , n12826 , n12832 , n12837 );
not ( n12839 , n12824 );
and ( n12840 , n12731 , n12839 , n987 );
nor ( n12841 , n1 , n12798 , n12746 );
nor ( n12842 , n12840 , n12841 );
not ( n12843 , n3609 );
not ( n12844 , n12823 );
or ( n12845 , n12843 , n12844 );
nand ( n12846 , n2506 , n12804 );
nand ( n12847 , n12845 , n12846 );
and ( n12848 , n12847 , n2298 , n12762 );
and ( n12849 , n2885 , n2508 , n5 , n12814 );
nor ( n12850 , n12848 , n12849 );
nand ( n12851 , n12819 , n12838 , n12842 , n12850 );
and ( n12852 , n3569 , n12851 );
or ( n12853 , n5 , n4183 );
nand ( n12854 , n2506 , n3754 );
nand ( n12855 , n12853 , n12854 );
and ( n12856 , n12855 , n12779 );
nor ( n12857 , n12852 , n12856 );
and ( n12858 , n12782 , n12789 , n12791 , n12857 );
nor ( n12859 , n7 , n12858 );
and ( n12860 , n4234 , n12859 );
nand ( n12861 , n10 , n4234 );
not ( n12862 , n12861 );
not ( n12863 , n3751 );
or ( n12864 , n445 , n13 );
nand ( n12865 , n12864 , n3117 );
and ( n12866 , n5897 , n12865 );
not ( n12867 , n2 );
not ( n12868 , n40 );
or ( n12869 , n12868 , n13 );
nand ( n12870 , n12869 , n1980 );
nand ( n12871 , n12867 , n12870 );
not ( n12872 , n2 );
nand ( n12873 , n12872 , n2308 );
and ( n12874 , n11 , n3914 );
nor ( n12875 , n12874 , n2 );
not ( n12876 , n12875 );
and ( n12877 , n12871 , n12873 , n12876 );
not ( n12878 , n12877 );
nand ( n12879 , n12866 , n12878 );
not ( n12880 , n2 );
not ( n12881 , n12880 );
not ( n12882 , n12708 );
or ( n12883 , n12881 , n12882 );
nand ( n12884 , n12883 , n12877 );
nand ( n12885 , n3609 , n12884 );
not ( n12886 , n986 );
not ( n12887 , n12886 );
not ( n12888 , n12766 );
or ( n12889 , n12887 , n12888 );
nand ( n12890 , n445 , n80 , n12752 );
nand ( n12891 , n12889 , n12890 );
nand ( n12892 , n39 , n12891 );
nand ( n12893 , n12879 , n12885 , n12892 );
and ( n12894 , n12863 , n12893 );
and ( n12895 , n12702 , n5313 );
nor ( n12896 , n12895 , n12772 );
or ( n12897 , n12702 , n5312 );
not ( n12898 , n13 );
not ( n12899 , n85 );
and ( n12900 , n12898 , n12899 );
not ( n12901 , n2 );
nor ( n12902 , n12901 , n2308 );
nor ( n12903 , n12900 , n12902 );
nand ( n12904 , n12897 , n12903 );
nor ( n12905 , n12875 , n12904 );
nand ( n12906 , n12896 , n12905 );
and ( n12907 , n3 , n12906 );
nor ( n12908 , n12894 , n12907 );
nand ( n12909 , n3753 , n4015 , n4157 , n12893 );
not ( n12910 , n3755 );
nand ( n12911 , n12910 , n12893 , n12866 );
and ( n12912 , n12908 , n12909 , n12911 );
and ( n12913 , n4166 , n5901 , n12720 );
and ( n12914 , n4167 , n12784 );
nand ( n12915 , n1852 , n2310 , n5314 );
not ( n12916 , n12915 );
nor ( n12917 , n12914 , n4159 , n12916 );
nor ( n12918 , n12913 , n12917 );
nand ( n12919 , n3753 , n5901 , n12720 );
nand ( n12920 , n4166 , n2508 , n4016 , n12915 );
and ( n12921 , n12912 , n12918 , n12919 , n12920 );
not ( n12922 , n12728 );
and ( n12923 , n12922 , n12891 );
and ( n12924 , n4252 , n12906 );
and ( n12925 , n39 , n4166 );
nor ( n12926 , n12925 , n12727 );
and ( n12927 , n41 , n12752 , n6440 );
nor ( n12928 , n41 , n4159 , n5898 );
nor ( n12929 , n12927 , n12928 );
or ( n12930 , n12926 , n12929 );
nand ( n12931 , n4166 , n2508 , n1971 , n5899 );
nand ( n12932 , n12930 , n12931 );
nor ( n12933 , n12923 , n12924 , n12932 );
and ( n12934 , n12752 , n6630 , n3750 );
and ( n12935 , n12934 , n3857 , n3531 );
nor ( n12936 , n41 , n5900 , n6860 );
and ( n12937 , n12936 , n2 , n4166 );
nor ( n12938 , n12935 , n12937 );
or ( n12939 , n3609 , n3569 , n2731 );
nand ( n12940 , n12939 , n4151 );
not ( n12941 , n12893 );
or ( n12942 , n3763 , n12941 );
and ( n12943 , n4015 , n12891 );
and ( n12944 , n39 , n12884 );
nor ( n12945 , n12943 , n12944 );
nand ( n12946 , n12877 , n12885 , n12892 );
nand ( n12947 , n12866 , n12946 );
nand ( n12948 , n12942 , n12945 , n12947 );
and ( n12949 , n12940 , n12948 );
nand ( n12950 , n6251 , n12854 );
and ( n12951 , n12950 , n12906 );
nor ( n12952 , n12949 , n12951 );
and ( n12953 , n12938 , n12952 );
nand ( n12954 , n12921 , n12933 , n12953 );
or ( n12955 , n5315 , n12735 );
nand ( n12956 , n12955 , n8 , n8885 );
nand ( n12957 , n8 , n8886 , n12777 );
nand ( n12958 , n12956 , n12957 );
nand ( n12959 , n10 , n12958 );
not ( n12960 , n12959 );
nor ( n12961 , n12862 , n7 , n12954 , n12960 );
nor ( n12962 , n7 , n8 );
nand ( n12963 , n10 , n4235 , n12954 );
and ( n12964 , n10 , n12962 , n12959 , n12963 );
nor ( n12965 , n12860 , n12961 , n12964 );
not ( n12966 , n12954 );
and ( n12967 , n12962 , n12959 , n12966 );
nand ( n12968 , n12963 , n12689 , n12959 );
or ( n12969 , n12858 , n12968 );
nand ( n12970 , n12969 , n9014 );
nor ( n12971 , n12967 , n12970 );
not ( n12972 , n4234 );
not ( n12973 , n12968 );
and ( n12974 , n12972 , n12973 );
not ( n12975 , n12859 );
or ( n12976 , n12975 , n12960 , n12954 );
or ( n12977 , n12691 , n12962 );
nand ( n12978 , n12977 , n4234 );
nand ( n12979 , n12976 , n12978 );
nor ( n12980 , n12974 , n12979 );
nand ( n12981 , n12697 , n12965 , n12971 , n12980 );
nand ( n12982 , n12681 , n12981 );
nand ( n12983 , n7 , n4235 );
nor ( n12984 , n31 , n12983 , n12695 );
or ( n12985 , n12958 , n12975 );
nand ( n12986 , n7 , n5821 , n12694 );
nor ( n12987 , n12692 , n12861 , n12986 );
nor ( n12988 , n6 , n12987 );
nor ( n12989 , n7 , n12958 );
and ( n12990 , n8 , n12989 );
and ( n12991 , n998 , n4235 , n12861 );
nor ( n12992 , n12991 , n12684 );
not ( n12993 , n12992 );
and ( n12994 , n7 , n12993 );
nor ( n12995 , n12990 , n12994 );
nand ( n12996 , n12985 , n12988 , n12995 );
or ( n12997 , n12984 , n12996 );
or ( n12998 , n9014 , n4235 );
nand ( n12999 , n12997 , n12998 );
or ( n13000 , n9014 , n4236 );
and ( n13001 , n12859 , n12959 , n12963 );
and ( n13002 , n8 , n12683 , n12695 );
nor ( n13003 , n13001 , n13002 );
not ( n13004 , n23 );
and ( n13005 , n13004 , n4234 , n12691 );
nor ( n13006 , n13005 , n6 );
or ( n13007 , n10 , n12684 );
nand ( n13008 , n13007 , n12685 );
and ( n13009 , n7 , n13008 );
and ( n13010 , n4235 , n4236 );
nand ( n13011 , n4235 , n4234 );
nor ( n13012 , n12692 , n13011 , n12986 );
nor ( n13013 , n13009 , n13010 , n13012 );
nand ( n13014 , n13003 , n12968 , n13006 , n13013 );
nand ( n13015 , n13000 , n13014 );
not ( n13016 , n9244 );
not ( n13017 , n13016 );
not ( n13018 , n13017 );
nor ( n13019 , n23 , n349 );
not ( n13020 , n13019 );
or ( n13021 , n13018 , n13020 );
nand ( n13022 , n22 , n348 );
and ( n13023 , n36 , n37 );
nor ( n13024 , n36 , n37 );
nor ( n13025 , n13023 , n13024 );
or ( n13026 , n31 , n13022 , n13025 );
nand ( n13027 , n13026 , n23 );
nand ( n13028 , n13021 , n13027 );
buf ( n13029 , n10240 );
buf ( n13030 , n13029 );
not ( n13031 , n13030 );
not ( n13032 , n13031 );
not ( n13033 , n7450 );
or ( n13034 , n13032 , n13033 );
nand ( n13035 , n13034 , n30 );
not ( n13036 , n13035 );
not ( n13037 , n33 );
and ( n13038 , n30 , n4512 );
nand ( n13039 , n13037 , n13038 );
not ( n13040 , n13031 );
not ( n13041 , n7448 );
not ( n13042 , n13041 );
or ( n13043 , n13040 , n13042 );
nand ( n13044 , n13043 , n30 );
and ( n13045 , n13036 , n13039 , n13044 );
buf ( n13046 , n13030 );
nand ( n13047 , n30 , n36 );
not ( n13048 , n13047 );
nor ( n13049 , n37 , n13048 );
not ( n13050 , n13049 );
not ( n13051 , n37 );
not ( n13052 , n30 );
nor ( n13053 , n13052 , n36 );
nor ( n13054 , n13051 , n13053 );
not ( n13055 , n13054 );
nand ( n13056 , n13050 , n13055 );
nand ( n13057 , n13046 , n13056 );
not ( n13058 , n13057 );
nor ( n13059 , n13045 , n13058 );
and ( n13060 , n14 , n13028 , n13059 );
nand ( n13061 , n13017 , n7353 );
not ( n13062 , n13061 );
not ( n13063 , n23 );
not ( n13064 , n13017 );
nor ( n13065 , n13064 , n10280 );
nand ( n13066 , n13062 , n14 , n13063 , n13065 );
or ( n13067 , n25 , n1054 );
not ( n13068 , n14 );
not ( n13069 , n23 );
not ( n13070 , n26 );
nand ( n13071 , n13069 , n13070 );
nor ( n13072 , n25 , n13068 , n13071 );
nand ( n13073 , n13065 , n13067 , n13072 );
nand ( n13074 , n13066 , n13073 );
nor ( n13075 , n13060 , n13074 );
or ( n13076 , n7838 , n13029 );
nand ( n13077 , n13076 , n30 );
and ( n13078 , n7444 , n13077 );
nor ( n13079 , n13078 , n34 );
and ( n13080 , n13079 , n13067 , n13072 );
not ( n13081 , n13079 );
nor ( n13082 , n13061 , n13081 );
not ( n13083 , n23 );
and ( n13084 , n13082 , n14 , n13083 );
nor ( n13085 , n13080 , n13084 );
not ( n13086 , n7521 );
not ( n13087 , n13067 );
nor ( n13088 , n23 , n13086 , n13087 );
and ( n13089 , n13088 , n14 , n13059 );
not ( n13090 , n13025 );
not ( n13091 , n13022 );
nand ( n13092 , n13090 , n5816 , n13091 );
nand ( n13093 , n3573 , n13092 );
not ( n13094 , n13093 );
nor ( n13095 , n13089 , n13094 );
and ( n13096 , n13075 , n13085 , n13095 );
not ( n13097 , n19 );
and ( n13098 , n46 , n13097 );
not ( n13099 , n13098 );
nor ( n13100 , n13096 , n13099 );
and ( n13101 , n20 , n13100 );
and ( n13102 , n30 , n34 );
nor ( n13103 , n13102 , n13029 );
nor ( n13104 , n7312 , n13103 );
nand ( n13105 , n34 , n13104 );
not ( n13106 , n33 );
nand ( n13107 , n13046 , n13047 );
nand ( n13108 , n13105 , n13106 , n13107 );
not ( n13109 , n34 );
or ( n13110 , n13030 , n13053 );
nand ( n13111 , n13110 , n7335 );
and ( n13112 , n13109 , n13111 );
or ( n13113 , n391 , n7323 );
nand ( n13114 , n13113 , n7444 );
and ( n13115 , n34 , n13114 );
or ( n13116 , n37 , n13112 , n13115 );
not ( n13117 , n13046 );
and ( n13118 , n37 , n393 );
nor ( n13119 , n13118 , n13024 );
or ( n13120 , n13117 , n13119 , n13115 );
nand ( n13121 , n13116 , n13120 );
and ( n13122 , n13108 , n13121 );
not ( n13123 , n13019 );
nand ( n13124 , n13123 , n13027 );
not ( n13125 , n33 );
nand ( n13126 , n232 , n13125 , n13108 );
not ( n13127 , n13044 );
nand ( n13128 , n37 , n13035 , n13039 , n13127 );
nand ( n13129 , n13124 , n13126 , n13128 );
nor ( n13130 , n13122 , n13129 );
not ( n13131 , n46 );
nor ( n13132 , n13131 , n14 );
not ( n13133 , n13117 );
nand ( n13134 , n13133 , n13054 );
and ( n13135 , n13130 , n13132 , n13134 );
not ( n13136 , n23 );
not ( n13137 , n13104 );
and ( n13138 , n13136 , n13087 , n13137 );
nor ( n13139 , n13138 , n13094 );
or ( n13140 , n13131 , n13139 );
not ( n13141 , n23 );
and ( n13142 , n13141 , n349 );
nand ( n13143 , n13132 , n13067 , n13142 , n13112 );
nand ( n13144 , n13140 , n13143 );
nor ( n13145 , n13135 , n13144 );
not ( n13146 , n13039 );
not ( n13147 , n13046 );
nand ( n13148 , n13147 , n9747 );
nand ( n13149 , n30 , n13148 );
nor ( n13150 , n13146 , n13149 );
or ( n13151 , n13046 , n9747 );
nand ( n13152 , n13151 , n30 );
and ( n13153 , n13150 , n37 , n13152 );
and ( n13154 , n232 , n13081 );
and ( n13155 , n13133 , n13049 );
nor ( n13156 , n13154 , n13155 );
not ( n13157 , n13108 );
nor ( n13158 , n13156 , n13115 , n13157 );
nor ( n13159 , n13153 , n13158 );
not ( n13160 , n14 );
nor ( n13161 , n13160 , n13131 );
and ( n13162 , n13161 , n13134 );
nand ( n13163 , n13159 , n13162 , n13126 , n13124 );
nand ( n13164 , n34 , n46 , n13142 , n13137 );
nand ( n13165 , n13161 , n13067 , n13142 , n13079 );
nand ( n13166 , n13145 , n13163 , n13164 , n13165 );
and ( n13167 , n453 , n13166 );
not ( n13168 , n4851 );
nand ( n13169 , n37 , n13168 , n13057 );
not ( n13170 , n19 );
or ( n13171 , n13169 , n13170 , n20 );
nand ( n13172 , n37 , n169 , n13057 );
or ( n13173 , n625 , n13172 );
nand ( n13174 , n13171 , n13173 );
and ( n13175 , n13124 , n13174 );
nor ( n13176 , n13101 , n13167 , n13175 );
not ( n13177 , n13176 );
not ( n13178 , n624 );
nor ( n13179 , n37 , n13178 );
and ( n13180 , n13115 , n13179 , n13124 );
and ( n13181 , n13137 , n626 , n13142 );
nor ( n13182 , n13180 , n13181 );
nand ( n13183 , n13057 , n13124 );
not ( n13184 , n13016 );
nand ( n13185 , n13184 , n13142 );
nand ( n13186 , n13183 , n13185 , n13093 );
and ( n13187 , n13131 , n20 , n13186 );
and ( n13188 , n908 , n13186 );
nor ( n13189 , n13187 , n13188 );
nand ( n13190 , n34 , n13107 );
nand ( n13191 , n13131 , n13190 , n13057 );
or ( n13192 , n13191 , n20 , n37 );
or ( n13193 , n46 , n20 , n13172 );
nand ( n13194 , n13192 , n13193 );
and ( n13195 , n13124 , n13194 );
and ( n13196 , n626 , n13094 );
nor ( n13197 , n13195 , n13196 );
not ( n13198 , n13168 );
nor ( n13199 , n46 , n13198 , n13183 );
not ( n13200 , n20 );
and ( n13201 , n13199 , n37 , n13200 );
and ( n13202 , n13142 , n13067 , n13065 );
nor ( n13203 , n10280 , n13185 );
nor ( n13204 , n13202 , n13203 );
not ( n13205 , n13112 );
and ( n13206 , n13079 , n13039 , n13205 );
nor ( n13207 , n13206 , n13058 );
and ( n13208 , n13028 , n13207 );
and ( n13209 , n13019 , n13207 );
not ( n13210 , n33 );
or ( n13211 , n13210 , n25 , n13071 );
nand ( n13212 , n13211 , n13185 );
and ( n13213 , n13112 , n13212 );
nor ( n13214 , n13208 , n13209 , n13213 );
and ( n13215 , n13204 , n13214 );
nand ( n13216 , n2382 , n13098 );
nor ( n13217 , n13215 , n13216 );
nor ( n13218 , n13201 , n13217 );
nand ( n13219 , n13182 , n13189 , n13197 , n13218 );
not ( n13220 , n20 );
and ( n13221 , n13220 , n13131 , n13142 , n13137 );
or ( n13222 , n46 , n20 , n13093 );
not ( n13223 , n13124 );
and ( n13224 , n13057 , n13179 , n13190 );
not ( n13225 , n13115 );
nor ( n13226 , n20 , n13225 );
and ( n13227 , n13226 , n232 , n13131 );
nor ( n13228 , n13224 , n13227 );
or ( n13229 , n13223 , n13228 );
nand ( n13230 , n13222 , n13229 );
nor ( n13231 , n13177 , n13219 , n13221 , n13230 );
nor ( n13232 , n5819 , n1868 );
not ( n13233 , n13232 );
or ( n13234 , n2385 , n13233 );
nand ( n13235 , n13234 , n841 );
and ( n13236 , n6833 , n13152 );
and ( n13237 , n13236 , n103 , n13039 );
and ( n13238 , n13152 , n103 , n3299 );
nor ( n13239 , n13237 , n13238 );
not ( n13240 , n33 );
and ( n13241 , n13240 , n101 );
and ( n13242 , n2816 , n13241 , n13039 );
not ( n13243 , n19 );
and ( n13244 , n13243 , n3815 );
nor ( n13245 , n13242 , n13244 );
nand ( n13246 , n13035 , n1866 , n8044 );
nand ( n13247 , n1866 , n13039 , n6725 , n13035 );
nand ( n13248 , n13239 , n13245 , n13246 , n13247 );
and ( n13249 , n391 , n1864 , n1919 );
and ( n13250 , n20 , n3815 );
nor ( n13251 , n13249 , n13250 );
nand ( n13252 , n33 , n101 );
not ( n13253 , n13252 );
nand ( n13254 , n642 , n13253 , n14 , n13044 );
not ( n13255 , n20 );
nor ( n13256 , n13255 , n16 );
nand ( n13257 , n14 , n13044 , n13256 , n13241 );
not ( n13258 , n20 );
nor ( n13259 , n13258 , n102 );
nand ( n13260 , n13149 , n13259 , n8044 );
and ( n13261 , n13251 , n13254 , n13257 , n13260 );
and ( n13262 , n13044 , n13259 , n3299 );
not ( n13263 , n33 );
and ( n13264 , n13263 , n2067 );
and ( n13265 , n33 , n912 );
nor ( n13266 , n13264 , n13265 );
and ( n13267 , n13266 , n391 , n103 );
nor ( n13268 , n13262 , n13267 );
not ( n13269 , n643 );
not ( n13270 , n14 );
nand ( n13271 , n13269 , n13253 , n13270 , n13149 );
not ( n13272 , n14 );
nand ( n13273 , n13256 , n13241 , n13272 , n13149 );
nand ( n13274 , n13261 , n13268 , n13271 , n13273 );
nor ( n13275 , n13248 , n13274 );
and ( n13276 , n13235 , n13275 );
not ( n13277 , n13038 );
nor ( n13278 , n13035 , n12383 , n3815 );
not ( n13279 , n13278 );
or ( n13280 , n13277 , n13279 );
nand ( n13281 , n2384 , n1870 , n13038 );
nand ( n13282 , n13280 , n13281 );
and ( n13283 , n13282 , n13275 );
not ( n13284 , n20 );
nor ( n13285 , n31 , n13241 );
not ( n13286 , n13248 );
nand ( n13287 , n2385 , n13285 , n13252 , n13286 );
and ( n13288 , n13284 , n13287 );
nor ( n13289 , n13288 , n13274 );
nor ( n13290 , n13276 , n13283 , n13289 );
not ( n13291 , n13253 );
not ( n13292 , n13285 );
and ( n13293 , n13291 , n13292 );
nor ( n13294 , n13293 , n2384 );
not ( n13295 , n3246 );
nor ( n13296 , n13152 , n13295 , n3815 );
or ( n13297 , n13294 , n13296 );
nand ( n13298 , n13297 , n13038 , n13275 );
or ( n13299 , n13296 , n13278 );
nand ( n13300 , n13299 , n13252 , n13275 );
nand ( n13301 , n13290 , n13298 , n13300 );
nand ( n13302 , n3 , n39 );
not ( n13303 , n13302 );
nand ( n13304 , n13303 , n34 , n12802 );
not ( n13305 , n298 );
nor ( n13306 , n13305 , n1864 );
or ( n13307 , n13304 , n2506 , n13306 );
nand ( n13308 , n24 , n22 , n34 );
or ( n13309 , n13308 , n4183 , n12802 );
nand ( n13310 , n13307 , n13309 );
and ( n13311 , n4266 , n13310 );
nand ( n13312 , n3 , n1866 );
not ( n13313 , n12802 );
nor ( n13314 , n39 , n13312 , n13313 );
and ( n13315 , n13314 , n1 , n34 );
nand ( n13316 , n998 , n102 );
not ( n13317 , n13316 );
nor ( n13318 , n4183 , n13317 );
and ( n13319 , n13318 , n34 , n13313 );
nor ( n13320 , n13315 , n13319 );
nand ( n13321 , n34 , n3908 , n4182 , n12802 );
nor ( n13322 , n8620 , n13313 );
nand ( n13323 , n1 , n3 , n34 , n13322 );
and ( n13324 , n13320 , n13321 , n13323 );
nor ( n13325 , n13324 , n4270 );
nand ( n13326 , n13306 , n12802 );
not ( n13327 , n13326 );
nor ( n13328 , n34 , n13327 );
nor ( n13329 , n40 , n13326 );
nor ( n13330 , n2298 , n1 );
and ( n13331 , n13330 , n4266 );
not ( n13332 , n4251 );
nand ( n13333 , n3 , n13332 );
and ( n13334 , n13333 , n4242 );
nor ( n13335 , n13331 , n13334 );
or ( n13336 , n13328 , n13329 , n13335 );
nand ( n13337 , n4266 , n3908 , n13317 );
or ( n13338 , n13337 , n4183 , n13313 );
nand ( n13339 , n13336 , n13338 );
nor ( n13340 , n13311 , n13325 , n13339 );
and ( n13341 , n34 , n4243 );
nor ( n13342 , n24 , n12802 );
not ( n13343 , n13342 );
nand ( n13344 , n1 , n4266 );
nor ( n13345 , n13343 , n13316 , n13344 , n13302 );
nor ( n13346 , n13341 , n13345 );
not ( n13347 , n24 );
not ( n13348 , n23 );
nor ( n13349 , n13348 , n31 );
nand ( n13350 , n13347 , n22 , n13349 );
nor ( n13351 , n13350 , n4270 );
nand ( n13352 , n39 , n12802 , n4182 , n13351 );
or ( n13353 , n6451 , n4270 , n4183 , n13326 );
nand ( n13354 , n13340 , n13346 , n13352 , n13353 );
not ( n13355 , n24 );
not ( n13356 , n22 );
and ( n13357 , n13356 , n8616 );
nand ( n13358 , n13355 , n13357 );
not ( n13359 , n35 );
and ( n13360 , n13358 , n13359 );
not ( n13361 , n13358 );
and ( n13362 , n13361 , n3836 );
nor ( n13363 , n13360 , n13362 );
and ( n13364 , n1845 , n993 );
nand ( n13365 , n4182 , n9012 );
not ( n13366 , n13365 );
nand ( n13367 , n4237 , n13366 );
nor ( n13368 , n13364 , n13367 );
and ( n13369 , n13363 , n13368 );
not ( n13370 , n22 );
and ( n13371 , n13370 , n13349 );
and ( n13372 , n41 , n13371 );
nand ( n13373 , n35 , n41 );
not ( n13374 , n13373 );
nor ( n13375 , n13372 , n13374 );
not ( n13376 , n13375 );
not ( n13377 , n13367 );
nand ( n13378 , n38 , n13376 , n12802 , n13377 );
not ( n13379 , n13 );
nand ( n13380 , n12 , n13379 );
nor ( n13381 , n3520 , n13380 , n13367 );
and ( n13382 , n13363 , n13381 );
and ( n13383 , n4182 , n4252 );
nand ( n13384 , n10074 , n4242 , n13375 );
nor ( n13385 , n13383 , n13313 , n13384 );
nor ( n13386 , n13382 , n13385 );
nand ( n13387 , n13378 , n13386 );
nor ( n13388 , n445 , n7919 );
nand ( n13389 , n38 , n41 );
nand ( n13390 , n13388 , n13389 , n13377 );
not ( n13391 , n12717 );
not ( n13392 , n13391 );
or ( n13393 , n13390 , n13392 , n13313 );
not ( n13394 , n35 );
or ( n13395 , n13394 , n4242 );
nand ( n13396 , n13393 , n13395 );
nor ( n13397 , n13369 , n13387 , n13396 );
not ( n13398 , n13388 );
nor ( n13399 , n13398 , n3819 , n4243 , n13366 );
and ( n13400 , n13399 , n5351 , n12802 );
not ( n13401 , n22 );
not ( n13402 , n13349 );
nor ( n13403 , n13401 , n13402 , n13367 );
nand ( n13404 , n35 , n13389 );
not ( n13405 , n13404 );
and ( n13406 , n13403 , n13405 , n12802 );
nor ( n13407 , n13400 , n13406 );
nand ( n13408 , n35 , n3820 , n13375 , n13365 );
not ( n13409 , n22 );
nand ( n13410 , n13409 , n13391 , n13389 , n12802 );
or ( n13411 , n13410 , n3836 , n24 );
or ( n13412 , n13404 , n13349 , n13313 );
nand ( n13413 , n13411 , n13412 );
and ( n13414 , n13377 , n13413 );
not ( n13415 , n35 );
or ( n13416 , n13415 , n12802 );
nand ( n13417 , n13416 , n13373 );
and ( n13418 , n13365 , n13417 );
nor ( n13419 , n13414 , n13418 );
nand ( n13420 , n13397 , n13407 , n13408 , n13419 );
and ( n13421 , n13358 , n32 );
not ( n13422 , n13358 );
and ( n13423 , n13422 , n39 );
nor ( n13424 , n13421 , n13423 );
not ( n13425 , n13424 );
and ( n13426 , n13425 , n13368 );
and ( n13427 , n32 , n4243 );
nor ( n13428 , n13426 , n13427 );
nor ( n13429 , n13367 , n13402 , n6451 );
and ( n13430 , n13429 , n7918 , n12802 );
not ( n13431 , n8621 );
nand ( n13432 , n32 , n13431 , n12802 );
nand ( n13433 , n39 , n40 , n12802 , n13357 );
and ( n13434 , n13432 , n13433 );
nor ( n13435 , n13434 , n13367 );
nor ( n13436 , n13430 , n13435 );
nand ( n13437 , n8618 , n12802 );
not ( n13438 , n13437 );
nand ( n13439 , n13438 , n7918 );
and ( n13440 , n32 , n13365 , n13439 );
not ( n13441 , n13365 );
not ( n13442 , n40 );
nor ( n13443 , n13441 , n13442 , n13439 , n4243 );
nor ( n13444 , n13440 , n13443 );
and ( n13445 , n12802 , n9835 , n13377 );
not ( n13446 , n3908 );
nand ( n13447 , n13446 , n13371 , n13377 );
or ( n13448 , n13447 , n12793 , n13313 );
not ( n13449 , n13381 );
or ( n13450 , n13424 , n13449 );
nand ( n13451 , n13448 , n13450 );
nor ( n13452 , n13445 , n13451 );
nand ( n13453 , n13428 , n13436 , n13444 , n13452 );
not ( n13454 , n14 );
nand ( n13455 , n13454 , n13098 );
not ( n13456 , n13455 );
nor ( n13457 , n10433 , n13025 );
and ( n13458 , n13371 , n13457 );
not ( n13459 , n13458 );
not ( n13460 , n23 );
and ( n13461 , n26 , n13460 , n13457 );
not ( n13462 , n23 );
or ( n13463 , n13462 , n9848 , n13025 );
not ( n13464 , n23 );
nor ( n13465 , n13464 , n102 );
or ( n13466 , n10247 , n13465 );
nand ( n13467 , n13463 , n13466 );
nor ( n13468 , n13461 , n13467 );
nand ( n13469 , n13459 , n13468 );
and ( n13470 , n13456 , n13469 );
not ( n13471 , n9320 );
nor ( n13472 , n13471 , n4351 );
not ( n13473 , n13472 );
or ( n13474 , n25 , n256 , n13455 );
not ( n13475 , n32 );
or ( n13476 , n13475 , n18 );
nand ( n13477 , n13474 , n13476 );
not ( n13478 , n13477 );
or ( n13479 , n13473 , n13478 );
not ( n13480 , n22 );
nor ( n13481 , n13402 , n13456 );
nand ( n13482 , n13480 , n13481 , n18 , n13457 );
nand ( n13483 , n13479 , n13482 );
nor ( n13484 , n13098 , n13468 );
nor ( n13485 , n13470 , n13483 , n13484 );
and ( n13486 , n13099 , n13458 );
not ( n13487 , n18 );
nor ( n13488 , n13487 , n13456 , n13468 );
nand ( n13489 , n35 , n9320 );
not ( n13490 , n13489 );
nand ( n13491 , n18 , n25 );
not ( n13492 , n13491 );
not ( n13493 , n9855 );
nand ( n13494 , n13490 , n13492 , n13493 , n13098 );
not ( n13495 , n14 );
nor ( n13496 , n13494 , n13495 , n26 );
nor ( n13497 , n13486 , n13488 , n13496 );
not ( n13498 , n10720 );
nand ( n13499 , n35 , n13472 , n13498 , n13456 );
not ( n13500 , n18 );
and ( n13501 , n13500 , n13098 , n13469 );
nor ( n13502 , n9855 , n13099 , n7439 );
not ( n13503 , n14 );
nor ( n13504 , n13503 , n18 );
and ( n13505 , n13502 , n13504 , n13472 );
nor ( n13506 , n13501 , n13505 );
nand ( n13507 , n13485 , n13497 , n13499 , n13506 );
and ( n13508 , n9037 , n294 );
not ( n13509 , n13357 );
nor ( n13510 , n13508 , n13509 );
or ( n13511 , n4334 , n9661 );
nand ( n13512 , n13511 , n25 );
nand ( n13513 , n18 , n22 );
or ( n13514 , n13512 , n13513 , n11429 );
not ( n13515 , n18 );
nand ( n13516 , n25 , n13515 , n1373 );
or ( n13517 , n32 , n13471 , n13516 );
nand ( n13518 , n13514 , n13517 );
not ( n13519 , n8044 );
or ( n13520 , n10454 , n13513 , n13519 );
not ( n13521 , n35 );
not ( n13522 , n22 );
nand ( n13523 , n13522 , n5817 );
nand ( n13524 , n13521 , n13523 );
or ( n13525 , n13491 , n2815 , n13524 );
nand ( n13526 , n13520 , n13525 );
nand ( n13527 , n18 , n5818 );
or ( n13528 , n11429 , n13527 , n13512 );
or ( n13529 , n13519 , n13527 , n10454 );
nand ( n13530 , n13528 , n13529 );
nor ( n13531 , n13510 , n13518 , n13526 , n13530 );
not ( n13532 , n18 );
nand ( n13533 , n13532 , n1373 , n13371 );
or ( n13534 , n9037 , n12383 , n13524 , n10454 );
nand ( n13535 , n35 , n13523 );
not ( n13536 , n13535 );
not ( n13537 , n14 );
nand ( n13538 , n13536 , n13537 , n9832 , n1554 );
not ( n13539 , n14 );
or ( n13540 , n13539 , n13512 , n294 , n13535 );
nand ( n13541 , n13533 , n13534 , n13538 , n13540 );
not ( n13542 , n22 );
or ( n13543 , n13542 , n1372 , n13491 );
nand ( n13544 , n1104 , n9320 );
or ( n13545 , n13544 , n13516 );
nand ( n13546 , n13543 , n13545 );
not ( n13547 , n13524 );
nand ( n13548 , n13547 , n19 , n9410 );
or ( n13549 , n13548 , n16 , n13512 );
or ( n13550 , n234 , n9037 , n13535 );
nand ( n13551 , n13549 , n13550 );
nor ( n13552 , n13541 , n13546 , n13551 );
not ( n13553 , n11086 );
nor ( n13554 , n35 , n13471 , n13553 );
not ( n13555 , n18 );
not ( n13556 , n26 );
and ( n13557 , n13556 , n465 );
nor ( n13558 , n13557 , n234 );
and ( n13559 , n13554 , n13555 , n13558 );
and ( n13560 , n1373 , n5820 , n13492 );
nor ( n13561 , n13559 , n13560 );
not ( n13562 , n18 );
and ( n13563 , n6835 , n13558 );
and ( n13564 , n11721 , n13493 );
nor ( n13565 , n13563 , n13564 );
or ( n13566 , n13489 , n13565 );
and ( n13567 , n3299 , n13558 );
and ( n13568 , n8044 , n13493 );
nor ( n13569 , n13567 , n13568 );
or ( n13570 , n13471 , n13569 );
and ( n13571 , n2332 , n13371 );
not ( n13572 , n9449 );
and ( n13573 , n25 , n9320 , n13572 );
nor ( n13574 , n13573 , n13371 );
or ( n13575 , n2815 , n13574 );
or ( n13576 , n234 , n35 , n2815 , n13544 );
nand ( n13577 , n13575 , n13576 );
nor ( n13578 , n13571 , n13577 );
nand ( n13579 , n13566 , n13570 , n13578 );
and ( n13580 , n13562 , n13579 );
not ( n13581 , n13493 );
not ( n13582 , n18 );
nor ( n13583 , n14 , n2384 );
nand ( n13584 , n13582 , n13583 );
nor ( n13585 , n13581 , n13471 , n13584 , n35 );
not ( n13586 , n32 );
and ( n13587 , n13586 , n25 , n10074 );
nor ( n13588 , n13587 , n13371 );
not ( n13589 , n32 );
and ( n13590 , n13589 , n25 , n1476 );
not ( n13591 , n32 );
nor ( n13592 , n13591 , n4367 , n13489 );
nor ( n13593 , n13590 , n13592 );
and ( n13594 , n13588 , n13593 );
not ( n13595 , n18 );
and ( n13596 , n13595 , n13583 );
and ( n13597 , n2385 , n13504 );
nor ( n13598 , n13596 , n13597 );
nor ( n13599 , n13594 , n13598 );
nor ( n13600 , n13580 , n13585 , n13599 );
nand ( n13601 , n13531 , n13552 , n13561 , n13600 );
and ( n13602 , n33 , n13437 );
and ( n13603 , n33 , n3819 );
nor ( n13604 , n13602 , n13603 );
not ( n13605 , n22 );
or ( n13606 , n13605 , n41 );
nand ( n13607 , n13606 , n33 );
nand ( n13608 , n41 , n12802 , n1869 , n5316 );
and ( n13609 , n13604 , n13607 , n13608 );
nor ( n13610 , n13609 , n13335 );
not ( n13611 , n13610 );
not ( n13612 , n22 );
nor ( n13613 , n23 , n24 );
or ( n13614 , n13612 , n13613 );
nand ( n13615 , n13614 , n33 );
or ( n13616 , n13615 , n4183 , n13313 );
not ( n13617 , n13312 );
nand ( n13618 , n41 , n13617 , n12802 );
not ( n13619 , n33 );
or ( n13620 , n13618 , n2506 , n13619 );
nand ( n13621 , n13616 , n13620 );
and ( n13622 , n4266 , n13621 );
nand ( n13623 , n33 , n13313 , n4182 , n13350 );
nand ( n13624 , n41 , n3836 , n4182 , n13327 );
and ( n13625 , n13623 , n13624 );
nor ( n13626 , n13625 , n4270 );
not ( n13627 , n13342 );
nand ( n13628 , n3 , n38 );
nor ( n13629 , n13627 , n13316 , n13344 , n13628 );
nor ( n13630 , n13622 , n13626 , n13629 );
and ( n13631 , n33 , n4243 );
nand ( n13632 , n12802 , n13351 );
or ( n13633 , n13632 , n2506 , n13628 );
nand ( n13634 , n4182 , n13316 , n12802 , n4266 );
not ( n13635 , n33 );
or ( n13636 , n13634 , n13635 , n38 );
nand ( n13637 , n13633 , n13636 );
not ( n13638 , n12802 );
not ( n13639 , n13389 );
not ( n13640 , n13316 );
and ( n13641 , n13639 , n13640 );
and ( n13642 , n33 , n13402 );
nor ( n13643 , n13641 , n13642 );
nor ( n13644 , n13638 , n4270 , n13643 , n4183 );
nor ( n13645 , n13631 , n13637 , n13644 );
nand ( n13646 , n13611 , n13630 , n13645 );
or ( n13647 , n1980 , n4230 );
or ( n13648 , n2 , n8841 );
nand ( n13649 , n40 , n11 , n12702 );
and ( n13650 , n2897 , n7794 );
not ( n13651 , n2 );
and ( n13652 , n13651 , n12801 );
nor ( n13653 , n13650 , n13652 );
nand ( n13654 , n13648 , n13649 , n13653 );
not ( n13655 , n13654 );
nand ( n13656 , n13655 , n4228 );
or ( n13657 , n2 , n13656 );
nand ( n13658 , n13 , n12682 );
nor ( n13659 , n12 , n6 , n13658 );
not ( n13660 , n13659 );
and ( n13661 , n12 , n2 , n1845 );
and ( n13662 , n2 , n4224 );
nor ( n13663 , n13661 , n13662 );
not ( n13664 , n13 );
or ( n13665 , n13664 , n3117 );
nand ( n13666 , n13665 , n2 );
nor ( n13667 , n1980 , n6 , n13658 );
and ( n13668 , n3796 , n13667 );
and ( n13669 , n3837 , n12902 );
nor ( n13670 , n13668 , n13669 );
nand ( n13671 , n13663 , n13666 , n13670 );
not ( n13672 , n13671 );
or ( n13673 , n13660 , n13672 );
nand ( n13674 , n13673 , n13380 );
nand ( n13675 , n12738 , n13649 , n13653 , n13674 );
nand ( n13676 , n13647 , n13657 , n13675 );
or ( n13677 , n2506 , n4230 );
and ( n13678 , n1 , n114 );
nor ( n13679 , n13678 , n5 );
or ( n13680 , n3609 , n4156 );
nand ( n13681 , n13680 , n6860 );
and ( n13682 , n4166 , n13681 );
or ( n13683 , n5 , n4182 );
nand ( n13684 , n5 , n4182 );
nand ( n13685 , n13683 , n13684 );
and ( n13686 , n3569 , n13685 );
nor ( n13687 , n13682 , n13686 );
or ( n13688 , n13679 , n13687 );
nor ( n13689 , n6855 , n13687 );
and ( n13690 , n2303 , n13689 );
nor ( n13691 , n2506 , n4 );
and ( n13692 , n13691 , n13687 );
nor ( n13693 , n13690 , n13692 );
nand ( n13694 , n4230 , n13688 , n2506 , n13693 );
nand ( n13695 , n13693 , n13691 , n13688 );
nand ( n13696 , n13677 , n13694 , n13695 );
not ( n13697 , n2 );
nor ( n13698 , n13697 , n4224 );
and ( n13699 , n2574 , n13698 );
and ( n13700 , n3523 , n13698 );
nand ( n13701 , n9 , n11666 );
or ( n13702 , n12684 , n13701 );
not ( n13703 , n13701 );
nand ( n13704 , n24 , n10431 );
nand ( n13705 , n13703 , n13704 , n13308 );
nand ( n13706 , n13702 , n13705 );
nor ( n13707 , n13700 , n13706 , n13667 );
and ( n13708 , n5817 , n13308 );
nor ( n13709 , n13708 , n9 );
not ( n13710 , n12983 );
and ( n13711 , n13709 , n9014 , n13710 );
not ( n13712 , n23 );
not ( n13713 , n8624 );
and ( n13714 , n13712 , n13713 );
nor ( n13715 , n13714 , n9 );
and ( n13716 , n13715 , n7 , n8 );
nor ( n13717 , n13711 , n13716 );
or ( n13718 , n10 , n5818 );
not ( n13719 , n13701 );
nand ( n13720 , n13718 , n13719 );
and ( n13721 , n11666 , n4237 );
and ( n13722 , n24 , n13704 );
or ( n13723 , n13722 , n11665 , n13011 );
or ( n13724 , n4235 , n11665 , n12861 );
nand ( n13725 , n13723 , n13724 );
nor ( n13726 , n13721 , n13725 , n6 );
nand ( n13727 , n13707 , n13717 , n13720 , n13726 );
not ( n13728 , n4226 );
nor ( n13729 , n13728 , n12877 );
nor ( n13730 , n13699 , n13727 , n13729 );
not ( n13731 , n3760 );
not ( n13732 , n2301 );
or ( n13733 , n13731 , n13732 );
nand ( n13734 , n13733 , n4 );
not ( n13735 , n13734 );
and ( n13736 , n13330 , n13735 );
nand ( n13737 , n4183 , n4226 , n114 , n6855 );
nor ( n13738 , n13737 , n4185 , n13734 );
nor ( n13739 , n1 , n6252 , n13735 );
nor ( n13740 , n13736 , n13738 , n13739 );
and ( n13741 , n3 , n4227 );
nand ( n13742 , n3569 , n114 , n13734 );
or ( n13743 , n13742 , n13728 , n4185 );
nor ( n13744 , n13330 , n4157 );
or ( n13745 , n13734 , n11376 , n13744 );
nand ( n13746 , n13743 , n13745 );
not ( n13747 , n13744 );
nand ( n13748 , n13747 , n3609 , n4249 );
or ( n13749 , n13748 , n2299 , n13734 );
not ( n13750 , n4167 );
nand ( n13751 , n13750 , n4183 , n4249 , n13734 );
nand ( n13752 , n13749 , n13751 );
nor ( n13753 , n13741 , n13746 , n13752 );
nand ( n13754 , n13740 , n13753 );
not ( n13755 , n13 );
not ( n13756 , n4229 );
or ( n13757 , n13755 , n13756 );
and ( n13758 , n13654 , n13659 , n12878 );
nor ( n13759 , n13 , n13728 , n13654 );
nor ( n13760 , n13758 , n13759 );
nor ( n13761 , n1845 , n12801 );
nand ( n13762 , n13654 , n13761 , n13729 );
nand ( n13763 , n13757 , n13760 , n13762 );
or ( n13764 , n1845 , n4228 );
or ( n13765 , n2 , n12878 );
not ( n13766 , n4225 );
nor ( n13767 , n11 , n3837 , n13766 );
or ( n13768 , n13761 , n13767 );
nand ( n13769 , n13765 , n13768 );
nand ( n13770 , n13764 , n13769 );
or ( n13771 , n3749 , n4183 , n4227 );
and ( n13772 , n13735 , n4226 , n13684 );
and ( n13773 , n4 , n4227 );
nor ( n13774 , n13772 , n13773 );
nand ( n13775 , n13771 , n13774 );
or ( n13776 , n7838 , n13232 );
nand ( n13777 , n13776 , n3821 );
nor ( n13778 , n3747 , n2898 , n4227 );
patch p0 (.w976043(t_0), .g0(g0), .g1(g1), .g2(g2), .g3(g3), .g4(g4), .g5(g5), .g6(g6), .g7(g7), .g8(g8), .g9(g9), .g10(g10), .g11(g11), .g12(g12), .g13(g13), .g14(g14), .g15(g15), .g16(g16), .g33(g33), .g17(g17), .g18(g18), .g19(g19), .g20(g20), .g21(g21), .g22(g22), .g23(g23), .g24(g24), .g25(g25), .g26(g26), .g27(g27), .g28(g28), .g29(g29), .g30(g30), .g31(g31), .g32(g32), .g34(g34), .g35(g35), .g36(g36), .g37(g37), .g38(g38), .g39(g39), .g40(g40), .g41(g41), .g42(g42), .g43(g43), .g44(g44), .g45(g45));
endmodule