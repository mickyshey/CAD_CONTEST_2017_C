module top (g32_po, g33_po, g34_po, g35_po, g36_po, g37_po, g38_po, g39_po, g40_po, g41_po, g42_po, g43_po, g44_po, g45_po, g46_po, g47_po, g48_po, g49_po, g50_po, g51_po, g52_po, g53_po, g54_po, g55_po, g56_po, g57_po, g58_po, g59_po, g60_po, g61_po, g62_po, g63_po, g64_po, g65_po, g66_po, g67_po, g68_po, g69_po, g70_po, g71_po, g72_po, g73_po, g74_po, g75_po, g76_po, g77_po, g78_po, g79_po, g80_po, g81_po, g82_po, g83_po, g84_po, g85_po, g86_po, g87_po, g88_po, g89_po, g90_po, g91_po, g92_po, g93_po, g94_po, g95_po, g96_po, g97_po, g98_po, g99_po, g100_po, g101_po, g102_po, g103_po, g104_po, g105_po, g106_po, g107_po, g108_po, g109_po, g110_po, g111_po, g112_po, g113_po, g114_po, g115_po, g116_po, g117_po, g118_po, g119_po, g120_po, g121_po, g122_po, g123_po, g124_po, g125_po, g126_po, g127_po, g128_po, g129_po, g130_po, g131_po, g132_po, g133_po, g134_po, g135_po, g136_po, g137_po, g138_po, g139_po, g140_po, g141_po, g142_po, g143_po, g144_po, g145_po, g146_po, g147_po, g148_po, g149_po, g150_po, g151_po, g152_po, g153_po, g154_po, g155_po, g156_po, g157_po, g158_po, g159_po, g160_po, g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g0_sel, g1_sel, g2_sel, g3_sel, g4_sel, g5_sel, g6_sel, g7_sel, g8_sel, g9_sel, g10_sel, g11_sel, g12_sel, g13_sel, g14_sel, g15_sel, g16_sel, g17_sel, g18_sel, g19_sel, g20_sel, g21_sel, g22_sel, g23_sel, g24_sel, g25_sel, g26_sel, g27_sel, g28_sel, g29_sel, g30_sel, g31_sel, g349_sel, g350_sel, g351_sel, g352_sel, g353_sel, g354_sel, g355_sel, g356_sel, g357_sel, n28_sel, n29_sel, n30_sel, n31_sel, n32_sel, n33_sel, n34_sel, n35_sel, n36_sel, n37_sel, n38_sel, n39_sel, n40_sel, n41_sel, n42_sel, n43_sel, n44_sel, n45_sel, n46_sel, n47_sel, n48_sel, n49_sel, n50_sel, n1349_sel, n966_sel, n592_sel, n1514_sel, n1132_sel, n747_sel, n378_sel, n1298_sel, n915_sel, n541_sel, g153_sel, n1464_sel, n1081_sel, n705_sel, n327_sel, n1247_sel, n27_sel, n490_sel, n1413_sel, n1030_sel, n654_sel, n1196_sel, n802_sel, n442_sel, n1362_sel, n979_sel, n605_sel, n1527_sel, n1145_sel, n12_sel, n391_sel, n1311_sel, n928_sel, n554_sel, n1476_sel, n1094_sel, n715_sel, n340_sel, n1260_sel, n877_sel, n503_sel, n1426_sel, n1043_sel, n667_sel, n1209_sel, n19_sel, n455_sel, n1375_sel, n992_sel, n618_sel, n1540_sel, n1158_sel, n770_sel, n404_sel, n1324_sel, n941_sel, n567_sel, n1489_sel, n1107_sel, n725_sel, n353_sel, n1273_sel, n890_sel, n516_sel, n1439_sel, n1056_sel, n680_sel, n302_sel, n1222_sel, n825_sel, n468_sel, n1388_sel, n1005_sel, n631_sel, n1553_sel, n1171_sel, n780_sel, n417_sel, n1337_sel, n954_sel, n580_sel, n1502_sel, n1120_sel, n738_sel, n366_sel, n1286_sel, n903_sel, n529_sel, n1452_sel, n1069_sel, n693_sel, n315_sel, n1235_sel, n835_sel, n478_sel, g90_sel, n1401_sel, n1018_sel, n642_sel, n1184_sel, n793_sel, n430_sel, n1350_sel, n967_sel, n593_sel, n1515_sel, n1133_sel, n748_sel, n379_sel, n1299_sel, n916_sel, n542_sel, g154_sel, n1465_sel, n1082_sel, n706_sel, n328_sel, n1248_sel, n845_sel, n491_sel, n1414_sel, n1031_sel, n655_sel, n1197_sel, n803_sel, n443_sel, n1363_sel, n980_sel, n606_sel, n1528_sel, n1146_sel, n758_sel, n392_sel, n1312_sel, n929_sel, n555_sel, n1477_sel, n1095_sel, n716_sel, n341_sel, n1261_sel, n878_sel, n504_sel, n1427_sel, n1044_sel, n668_sel, n1210_sel, n20_sel, n456_sel, n1376_sel, n993_sel, n619_sel, n1541_sel, n1159_sel, n771_sel, n405_sel, n1325_sel, n942_sel, n568_sel, n1490_sel, n1108_sel, n726_sel, n354_sel, n1274_sel, n891_sel, n517_sel, n1440_sel, n1057_sel, n681_sel, n303_sel, n1223_sel, n826_sel, n469_sel, n1389_sel, n1006_sel, n632_sel, n1554_sel, n1172_sel, n781_sel, n418_sel, n1338_sel, n955_sel, n581_sel, n1503_sel, n1121_sel, n7_sel, n367_sel, n1287_sel, n904_sel, n530_sel, n1453_sel, n1070_sel, n694_sel, n316_sel, n1236_sel, n836_sel, n479_sel, g91_sel, n1402_sel, n1019_sel, n643_sel, n1185_sel, n794_sel, n431_sel, n1351_sel, n968_sel, n594_sel, n1516_sel, n1134_sel, n749_sel, n380_sel, n1300_sel, n917_sel, n543_sel, g155_sel, n1466_sel, n1083_sel, n1_sel, n329_sel, n1249_sel, n866_sel, n492_sel, n1415_sel, n1032_sel, n656_sel, n1198_sel, n444_sel, n804_sel, n1364_sel, n981_sel, n607_sel, n1529_sel, n1147_sel, n393_sel, n759_sel, n1313_sel, n930_sel, n556_sel, n1478_sel, n1096_sel, n717_sel, n342_sel, n1262_sel, n879_sel, n505_sel, n1428_sel, n1045_sel, n669_sel, n1211_sel, n21_sel, n457_sel, n1377_sel, n994_sel, n620_sel, n1542_sel, n1160_sel, n406_sel, n772_sel, n1326_sel, n943_sel, n569_sel, n1491_sel, n1109_sel, n355_sel, n727_sel, n1275_sel, n892_sel, n518_sel, n1441_sel, n1058_sel, n304_sel, n682_sel, n1224_sel, n827_sel, n470_sel, n1390_sel, n1007_sel, n633_sel, n1555_sel, n1173_sel, n419_sel, n782_sel, n1339_sel, n956_sel, n582_sel, n1504_sel, n1122_sel, n368_sel, n8_sel, n1288_sel, n905_sel, n531_sel, n1454_sel, n1071_sel, n317_sel, n695_sel, n1237_sel, n837_sel, n480_sel, g92_sel, n1403_sel, n1020_sel, n644_sel, n1186_sel, n432_sel, n795_sel, n1352_sel, n969_sel, n595_sel, n1517_sel, n1135_sel, n381_sel, n750_sel, n1301_sel, n918_sel, g156_sel, n544_sel, n1467_sel, n1084_sel, n330_sel, n2_sel, n1250_sel, n867_sel, n493_sel, n1416_sel, n1033_sel, n657_sel, n1199_sel, n805_sel, n445_sel, n1365_sel, n982_sel, n608_sel, n1530_sel, n1148_sel, n760_sel, n394_sel, n1314_sel, n931_sel, n557_sel, n1479_sel, n1097_sel, n343_sel, n718_sel, n1263_sel, n880_sel, n506_sel, n1429_sel, n1046_sel, n670_sel, n1212_sel, n815_sel, n458_sel, n1378_sel, n995_sel, n621_sel, n1543_sel, n1161_sel, n773_sel, n407_sel, n1327_sel, n944_sel, n570_sel, n1492_sel, n1110_sel, n728_sel, n356_sel, n1276_sel, n893_sel, n519_sel, n1442_sel, n1059_sel, n683_sel, n305_sel, n1225_sel, n828_sel, g80_sel, n1391_sel, n1008_sel, n634_sel, n1556_sel, n1174_sel, n783_sel, n420_sel, n1340_sel, n957_sel, n583_sel, n1505_sel, n1123_sel, n9_sel, n369_sel, n1289_sel, n906_sel, g144_sel, n532_sel, n1455_sel, n1072_sel, n696_sel, n318_sel, n1238_sel, n838_sel, g93_sel, n481_sel, n1404_sel, n1021_sel, n645_sel, n1187_sel, n16_sel, n433_sel, n1353_sel, n970_sel, n596_sel, n1518_sel, n1136_sel, n751_sel, n382_sel, n1302_sel, n919_sel, n545_sel, g157_sel, n1468_sel, n1085_sel, n3_sel, n331_sel, n1251_sel, n868_sel, n494_sel, n1417_sel, n1034_sel, n658_sel, n1200_sel, n806_sel, n446_sel, n1366_sel, n983_sel, n609_sel, n1531_sel, n1149_sel, n761_sel, n395_sel, n1315_sel, n932_sel, n558_sel, n1480_sel, n1098_sel, n719_sel, n344_sel, n1264_sel, n881_sel, n507_sel, n1430_sel, n1047_sel, n671_sel, n1213_sel, n816_sel, n459_sel, n1379_sel, n996_sel, n622_sel, n1544_sel, n1162_sel, n774_sel, n408_sel, n1328_sel, n945_sel, n571_sel, n1493_sel, n1111_sel, n729_sel, n357_sel, n1277_sel, n894_sel, n520_sel, n1443_sel, n1060_sel, n684_sel, n306_sel, n1226_sel, n829_sel, g81_sel, n1392_sel, n1009_sel, n635_sel, n1557_sel, n1175_sel, n784_sel, n421_sel, n1341_sel, n958_sel, n584_sel, n1506_sel, n1124_sel, n739_sel, n370_sel, n1290_sel, n907_sel, n533_sel, g145_sel, n1456_sel, n1073_sel, n697_sel, n319_sel, n1239_sel, n839_sel, n482_sel, g94_sel, n1405_sel, n1022_sel, n646_sel, n1188_sel, n17_sel, n434_sel, n1354_sel, n971_sel, n597_sel, n1519_sel, n1137_sel, n752_sel, n383_sel, n1303_sel, n920_sel, n546_sel, g158_sel, n1469_sel, n1086_sel, n707_sel, n332_sel, n1252_sel, n869_sel, n495_sel, n1418_sel, n1035_sel, n659_sel, n1201_sel, n807_sel, n447_sel, n1367_sel, n984_sel, n610_sel, n1532_sel, n1150_sel, n762_sel, n396_sel, n1316_sel, n933_sel, n559_sel, n1481_sel, n1099_sel, n4_sel, n345_sel, n1265_sel, n882_sel, n508_sel, n1431_sel, n1048_sel, n672_sel, n1214_sel, n817_sel, n460_sel, n1380_sel, n997_sel, n623_sel, n1545_sel, n1163_sel, n775_sel, n409_sel, n1329_sel, n946_sel, n572_sel, n1494_sel, n1112_sel, n730_sel, n358_sel, n1278_sel, n895_sel, n521_sel, n1444_sel, n1061_sel, n685_sel, n307_sel, n1227_sel, n830_sel, g82_sel, n1393_sel, n1010_sel, n636_sel, n1558_sel, n1176_sel, n785_sel, n422_sel, n1342_sel, n959_sel, n585_sel, n1507_sel, n1125_sel, n740_sel, n371_sel, n1291_sel, n908_sel, n534_sel, g146_sel, n1457_sel, n1074_sel, n698_sel, n320_sel, n1240_sel, n840_sel, n483_sel, g95_sel, n1406_sel, n1023_sel, n647_sel, n1189_sel, n18_sel, n435_sel, n1355_sel, n972_sel, n598_sel, n1520_sel, n1138_sel, n753_sel, n384_sel, n1304_sel, n921_sel, n547_sel, g159_sel, n1470_sel, n1087_sel, n708_sel, n333_sel, n1253_sel, n870_sel, n496_sel, n1419_sel, n1036_sel, n660_sel, n1202_sel, n808_sel, n448_sel, n1368_sel, n985_sel, n611_sel, n1533_sel, n1151_sel, n763_sel, n397_sel, n1317_sel, n934_sel, n560_sel, n1482_sel, n1100_sel, n5_sel, n346_sel, n1266_sel, n883_sel, n509_sel, n1432_sel, n1049_sel, n673_sel, n1215_sel, n818_sel, n461_sel, n1381_sel, n998_sel, n624_sel, n1546_sel, n1164_sel, n776_sel, n410_sel, n1330_sel, n947_sel, n573_sel, n1495_sel, n1113_sel, n731_sel, n359_sel, n1279_sel, n896_sel, n522_sel, n1445_sel, n1062_sel, n686_sel, n308_sel, n1228_sel, n831_sel, n471_sel, g83_sel, n1394_sel, n1011_sel, n637_sel, n1177_sel, n786_sel, n423_sel, n1343_sel, n960_sel, n586_sel, n1508_sel, n1126_sel, n741_sel, n372_sel, n1292_sel, n909_sel, n535_sel, g147_sel, n1458_sel, n1075_sel, n699_sel, n321_sel, n1241_sel, n841_sel, n484_sel, g96_sel, n1407_sel, n1024_sel, n648_sel, n1190_sel, n796_sel, n436_sel, n1356_sel, n973_sel, n599_sel, n1521_sel, n1139_sel, n754_sel, n385_sel, n1305_sel, n922_sel, n548_sel, g160_sel, n1088_sel, n709_sel, n334_sel, n1254_sel, n871_sel, n497_sel, n1420_sel, n1037_sel, n661_sel, n1203_sel, n809_sel, n449_sel, n1369_sel, n986_sel, n612_sel, n1534_sel, n1152_sel, n764_sel, n398_sel, n1318_sel, n935_sel, n561_sel, n1483_sel, n1101_sel, n6_sel, n347_sel, n1267_sel, n884_sel, n510_sel, n1433_sel, n1050_sel, n674_sel, n1216_sel, n819_sel, n462_sel, n1382_sel, n999_sel, n625_sel, n1547_sel, n1165_sel, n13_sel, n411_sel, n1331_sel, n948_sel, n574_sel, n1496_sel, n1114_sel, n732_sel, n360_sel, n1280_sel, n897_sel, n523_sel, n1446_sel, n1063_sel, n687_sel, n309_sel, n1229_sel, n832_sel, n472_sel, g84_sel, n1395_sel, n1012_sel, n1178_sel, n787_sel, n424_sel, n1344_sel, n961_sel, n587_sel, n1509_sel, n1127_sel, n742_sel, n373_sel, n1293_sel, n910_sel, n536_sel, g148_sel, n1459_sel, n1076_sel, n700_sel, n322_sel, n1242_sel, n842_sel, n485_sel, n1408_sel, n1025_sel, n649_sel, n1191_sel, n797_sel, n437_sel, n1357_sel, n974_sel, n600_sel, n1522_sel, n1140_sel, n755_sel, n386_sel, n1306_sel, n923_sel, n549_sel, n1471_sel, n1089_sel, n710_sel, n335_sel, n1255_sel, n872_sel, n498_sel, n1421_sel, n1038_sel, n662_sel, n1204_sel, n810_sel, n450_sel, n1370_sel, n987_sel, n613_sel, n1535_sel, n1153_sel, n765_sel, n399_sel, n1319_sel, n936_sel, n562_sel, n1484_sel, n1102_sel, n720_sel, n348_sel, n1268_sel, n885_sel, n511_sel, n1434_sel, n1051_sel, n675_sel, n1217_sel, n820_sel, n463_sel, n1383_sel, n1000_sel, n626_sel, n1548_sel, n1166_sel, n14_sel, n412_sel, n1332_sel, n949_sel, n575_sel, n1497_sel, n1115_sel, n733_sel, n361_sel, n1281_sel, n898_sel, n524_sel, n1447_sel, n1064_sel, n688_sel, n310_sel, n1230_sel, n833_sel, n473_sel, g85_sel, n1396_sel, n1013_sel, n1179_sel, n425_sel, n788_sel, n1345_sel, n962_sel, n588_sel, n1510_sel, n1128_sel, n374_sel, n743_sel, n1294_sel, n911_sel, n537_sel, g149_sel, n1460_sel, n1077_sel, n323_sel, n701_sel, n1243_sel, n843_sel, n486_sel, n1409_sel, n1026_sel, n650_sel, n1192_sel, n438_sel, n798_sel, n1358_sel, n975_sel, n601_sel, n1523_sel, n1141_sel, n387_sel, n756_sel, n1307_sel, n924_sel, n550_sel, n1472_sel, n1090_sel, n336_sel, n711_sel, n1256_sel, n873_sel, n499_sel, n1422_sel, n1039_sel, n663_sel, n1205_sel, n451_sel, n811_sel, n1371_sel, n988_sel, n614_sel, n1536_sel, n1154_sel, n400_sel, n766_sel, n1320_sel, n937_sel, n563_sel, n1485_sel, n1103_sel, n349_sel, n721_sel, n1269_sel, n886_sel, n512_sel, n1435_sel, n1052_sel, n298_sel, n676_sel, n1218_sel, n821_sel, n464_sel, n1384_sel, n1001_sel, n627_sel, n1549_sel, n1167_sel, n413_sel, n15_sel, n1333_sel, n950_sel, n576_sel, n1498_sel, n1116_sel, n362_sel, n734_sel, n1282_sel, n899_sel, n525_sel, n1448_sel, n1065_sel, n311_sel, n689_sel, n1231_sel, n22_sel, g86_sel, n474_sel, n1397_sel, n1014_sel, n638_sel, n1180_sel, n789_sel, n426_sel, n1346_sel, n963_sel, n589_sel, n1511_sel, n1129_sel, n744_sel, n375_sel, n1295_sel, n912_sel, g150_sel, n538_sel, n1461_sel, n1078_sel, n702_sel, n324_sel, n1244_sel, n844_sel, n487_sel, n1410_sel, n1027_sel, n651_sel, n1193_sel, n799_sel, n439_sel, n1359_sel, n976_sel, n602_sel, n1524_sel, n1142_sel, n757_sel, n388_sel, n1308_sel, n925_sel, n551_sel, n1473_sel, n1091_sel, n712_sel, n337_sel, n1257_sel, n874_sel, n500_sel, n1423_sel, n1040_sel, n664_sel, n1206_sel, n812_sel, n452_sel, n1372_sel, n989_sel, n615_sel, n1537_sel, n1155_sel, n767_sel, n401_sel, n1321_sel, n938_sel, n564_sel, n1486_sel, n1104_sel, n722_sel, n350_sel, n1270_sel, n887_sel, n513_sel, n1436_sel, n1053_sel, n677_sel, n299_sel, n1219_sel, n822_sel, n465_sel, n1385_sel, n1002_sel, n628_sel, n1550_sel, n1168_sel, n777_sel, n414_sel, n1334_sel, n951_sel, n577_sel, n1499_sel, n1117_sel, n735_sel, n363_sel, n1283_sel, n900_sel, n526_sel, n1449_sel, n1066_sel, n690_sel, n312_sel, n1232_sel, n23_sel, n475_sel, g87_sel, n1398_sel, n1015_sel, n639_sel, n1181_sel, n790_sel, n427_sel, n1347_sel, n964_sel, n590_sel, n1512_sel, n1130_sel, n745_sel, n376_sel, n1296_sel, n913_sel, n539_sel, g151_sel, n1462_sel, n1079_sel, n703_sel, n325_sel, n1245_sel, n25_sel, n488_sel, n1411_sel, n1028_sel, n652_sel, n1194_sel, n800_sel, n440_sel, n1360_sel, n977_sel, n603_sel, n1525_sel, n1143_sel, n10_sel, n389_sel, n1309_sel, n926_sel, n552_sel, n1474_sel, n1092_sel, n713_sel, n338_sel, n1258_sel, n875_sel, n501_sel, n1424_sel, n1041_sel, n665_sel, n1207_sel, n813_sel, n453_sel, n1373_sel, n990_sel, n616_sel, n1538_sel, n1156_sel, n768_sel, n402_sel, n1322_sel, n939_sel, n565_sel, n1487_sel, n1105_sel, n723_sel, n351_sel, n1271_sel, n888_sel, n514_sel, n1437_sel, n1054_sel, n678_sel, n300_sel, n1220_sel, n823_sel, n466_sel, n1386_sel, n1003_sel, n629_sel, n1551_sel, n1169_sel, n778_sel, n415_sel, n1335_sel, n952_sel, n578_sel, n1500_sel, n1118_sel, n736_sel, n364_sel, n1284_sel, n901_sel, n527_sel, n1450_sel, n1067_sel, n691_sel, n313_sel, n1233_sel, n24_sel, n476_sel, g88_sel, n1399_sel, n1016_sel, n640_sel, n1182_sel, n791_sel, n428_sel, n1348_sel, n965_sel, n591_sel, n1513_sel, n1131_sel, n746_sel, n377_sel, n1297_sel, n914_sel, n540_sel, g152_sel, n1463_sel, n1080_sel, n704_sel, n326_sel, n1246_sel, n26_sel, n489_sel, n1412_sel, n1029_sel, n653_sel, n1195_sel, n801_sel, n441_sel, n1361_sel, n978_sel, n604_sel, n1526_sel, n1144_sel, n11_sel, n390_sel, n1310_sel, n927_sel, n553_sel, n1475_sel, n1093_sel, n714_sel, n339_sel, n1259_sel, n876_sel, n502_sel, n1425_sel, n1042_sel, n666_sel, n1208_sel, n814_sel, n454_sel, n1374_sel, n991_sel, n617_sel, n1539_sel, n1157_sel, n769_sel, n403_sel, n1323_sel, n940_sel, n566_sel, n1488_sel, n1106_sel, n724_sel, n352_sel, n1272_sel, n889_sel, n515_sel, n1438_sel, n1055_sel, n679_sel, n301_sel, n1221_sel, n824_sel, n467_sel, n1387_sel, n1004_sel, n630_sel, n1552_sel, n1170_sel, n779_sel, n416_sel, n1336_sel, n953_sel, n579_sel, n1501_sel, n1119_sel, n737_sel, n365_sel, n1285_sel, n902_sel, n528_sel, n1451_sel, n1068_sel, n692_sel, n314_sel, n1234_sel, n834_sel, n477_sel, g89_sel, n1400_sel, n1017_sel, n641_sel, n1183_sel, n792_sel, n429_sel);
input g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g0_sel, g1_sel, g2_sel, g3_sel, g4_sel, g5_sel, g6_sel, g7_sel, g8_sel, g9_sel, g10_sel, g11_sel, g12_sel, g13_sel, g14_sel, g15_sel, g16_sel, g17_sel, g18_sel, g19_sel, g20_sel, g21_sel, g22_sel, g23_sel, g24_sel, g25_sel, g26_sel, g27_sel, g28_sel, g29_sel, g30_sel, g31_sel, g349_sel, g350_sel, g351_sel, g352_sel, g353_sel, g354_sel, g355_sel, g356_sel, g357_sel, n28_sel, n29_sel, n30_sel, n31_sel, n32_sel, n33_sel, n34_sel, n35_sel, n36_sel, n37_sel, n38_sel, n39_sel, n40_sel, n41_sel, n42_sel, n43_sel, n44_sel, n45_sel, n46_sel, n47_sel, n48_sel, n49_sel, n50_sel, n1349_sel, n966_sel, n592_sel, n1514_sel, n1132_sel, n747_sel, n378_sel, n1298_sel, n915_sel, n541_sel, g153_sel, n1464_sel, n1081_sel, n705_sel, n327_sel, n1247_sel, n27_sel, n490_sel, n1413_sel, n1030_sel, n654_sel, n1196_sel, n802_sel, n442_sel, n1362_sel, n979_sel, n605_sel, n1527_sel, n1145_sel, n12_sel, n391_sel, n1311_sel, n928_sel, n554_sel, n1476_sel, n1094_sel, n715_sel, n340_sel, n1260_sel, n877_sel, n503_sel, n1426_sel, n1043_sel, n667_sel, n1209_sel, n19_sel, n455_sel, n1375_sel, n992_sel, n618_sel, n1540_sel, n1158_sel, n770_sel, n404_sel, n1324_sel, n941_sel, n567_sel, n1489_sel, n1107_sel, n725_sel, n353_sel, n1273_sel, n890_sel, n516_sel, n1439_sel, n1056_sel, n680_sel, n302_sel, n1222_sel, n825_sel, n468_sel, n1388_sel, n1005_sel, n631_sel, n1553_sel, n1171_sel, n780_sel, n417_sel, n1337_sel, n954_sel, n580_sel, n1502_sel, n1120_sel, n738_sel, n366_sel, n1286_sel, n903_sel, n529_sel, n1452_sel, n1069_sel, n693_sel, n315_sel, n1235_sel, n835_sel, n478_sel, g90_sel, n1401_sel, n1018_sel, n642_sel, n1184_sel, n793_sel, n430_sel, n1350_sel, n967_sel, n593_sel, n1515_sel, n1133_sel, n748_sel, n379_sel, n1299_sel, n916_sel, n542_sel, g154_sel, n1465_sel, n1082_sel, n706_sel, n328_sel, n1248_sel, n845_sel, n491_sel, n1414_sel, n1031_sel, n655_sel, n1197_sel, n803_sel, n443_sel, n1363_sel, n980_sel, n606_sel, n1528_sel, n1146_sel, n758_sel, n392_sel, n1312_sel, n929_sel, n555_sel, n1477_sel, n1095_sel, n716_sel, n341_sel, n1261_sel, n878_sel, n504_sel, n1427_sel, n1044_sel, n668_sel, n1210_sel, n20_sel, n456_sel, n1376_sel, n993_sel, n619_sel, n1541_sel, n1159_sel, n771_sel, n405_sel, n1325_sel, n942_sel, n568_sel, n1490_sel, n1108_sel, n726_sel, n354_sel, n1274_sel, n891_sel, n517_sel, n1440_sel, n1057_sel, n681_sel, n303_sel, n1223_sel, n826_sel, n469_sel, n1389_sel, n1006_sel, n632_sel, n1554_sel, n1172_sel, n781_sel, n418_sel, n1338_sel, n955_sel, n581_sel, n1503_sel, n1121_sel, n7_sel, n367_sel, n1287_sel, n904_sel, n530_sel, n1453_sel, n1070_sel, n694_sel, n316_sel, n1236_sel, n836_sel, n479_sel, g91_sel, n1402_sel, n1019_sel, n643_sel, n1185_sel, n794_sel, n431_sel, n1351_sel, n968_sel, n594_sel, n1516_sel, n1134_sel, n749_sel, n380_sel, n1300_sel, n917_sel, n543_sel, g155_sel, n1466_sel, n1083_sel, n1_sel, n329_sel, n1249_sel, n866_sel, n492_sel, n1415_sel, n1032_sel, n656_sel, n1198_sel, n444_sel, n804_sel, n1364_sel, n981_sel, n607_sel, n1529_sel, n1147_sel, n393_sel, n759_sel, n1313_sel, n930_sel, n556_sel, n1478_sel, n1096_sel, n717_sel, n342_sel, n1262_sel, n879_sel, n505_sel, n1428_sel, n1045_sel, n669_sel, n1211_sel, n21_sel, n457_sel, n1377_sel, n994_sel, n620_sel, n1542_sel, n1160_sel, n406_sel, n772_sel, n1326_sel, n943_sel, n569_sel, n1491_sel, n1109_sel, n355_sel, n727_sel, n1275_sel, n892_sel, n518_sel, n1441_sel, n1058_sel, n304_sel, n682_sel, n1224_sel, n827_sel, n470_sel, n1390_sel, n1007_sel, n633_sel, n1555_sel, n1173_sel, n419_sel, n782_sel, n1339_sel, n956_sel, n582_sel, n1504_sel, n1122_sel, n368_sel, n8_sel, n1288_sel, n905_sel, n531_sel, n1454_sel, n1071_sel, n317_sel, n695_sel, n1237_sel, n837_sel, n480_sel, g92_sel, n1403_sel, n1020_sel, n644_sel, n1186_sel, n432_sel, n795_sel, n1352_sel, n969_sel, n595_sel, n1517_sel, n1135_sel, n381_sel, n750_sel, n1301_sel, n918_sel, g156_sel, n544_sel, n1467_sel, n1084_sel, n330_sel, n2_sel, n1250_sel, n867_sel, n493_sel, n1416_sel, n1033_sel, n657_sel, n1199_sel, n805_sel, n445_sel, n1365_sel, n982_sel, n608_sel, n1530_sel, n1148_sel, n760_sel, n394_sel, n1314_sel, n931_sel, n557_sel, n1479_sel, n1097_sel, n343_sel, n718_sel, n1263_sel, n880_sel, n506_sel, n1429_sel, n1046_sel, n670_sel, n1212_sel, n815_sel, n458_sel, n1378_sel, n995_sel, n621_sel, n1543_sel, n1161_sel, n773_sel, n407_sel, n1327_sel, n944_sel, n570_sel, n1492_sel, n1110_sel, n728_sel, n356_sel, n1276_sel, n893_sel, n519_sel, n1442_sel, n1059_sel, n683_sel, n305_sel, n1225_sel, n828_sel, g80_sel, n1391_sel, n1008_sel, n634_sel, n1556_sel, n1174_sel, n783_sel, n420_sel, n1340_sel, n957_sel, n583_sel, n1505_sel, n1123_sel, n9_sel, n369_sel, n1289_sel, n906_sel, g144_sel, n532_sel, n1455_sel, n1072_sel, n696_sel, n318_sel, n1238_sel, n838_sel, g93_sel, n481_sel, n1404_sel, n1021_sel, n645_sel, n1187_sel, n16_sel, n433_sel, n1353_sel, n970_sel, n596_sel, n1518_sel, n1136_sel, n751_sel, n382_sel, n1302_sel, n919_sel, n545_sel, g157_sel, n1468_sel, n1085_sel, n3_sel, n331_sel, n1251_sel, n868_sel, n494_sel, n1417_sel, n1034_sel, n658_sel, n1200_sel, n806_sel, n446_sel, n1366_sel, n983_sel, n609_sel, n1531_sel, n1149_sel, n761_sel, n395_sel, n1315_sel, n932_sel, n558_sel, n1480_sel, n1098_sel, n719_sel, n344_sel, n1264_sel, n881_sel, n507_sel, n1430_sel, n1047_sel, n671_sel, n1213_sel, n816_sel, n459_sel, n1379_sel, n996_sel, n622_sel, n1544_sel, n1162_sel, n774_sel, n408_sel, n1328_sel, n945_sel, n571_sel, n1493_sel, n1111_sel, n729_sel, n357_sel, n1277_sel, n894_sel, n520_sel, n1443_sel, n1060_sel, n684_sel, n306_sel, n1226_sel, n829_sel, g81_sel, n1392_sel, n1009_sel, n635_sel, n1557_sel, n1175_sel, n784_sel, n421_sel, n1341_sel, n958_sel, n584_sel, n1506_sel, n1124_sel, n739_sel, n370_sel, n1290_sel, n907_sel, n533_sel, g145_sel, n1456_sel, n1073_sel, n697_sel, n319_sel, n1239_sel, n839_sel, n482_sel, g94_sel, n1405_sel, n1022_sel, n646_sel, n1188_sel, n17_sel, n434_sel, n1354_sel, n971_sel, n597_sel, n1519_sel, n1137_sel, n752_sel, n383_sel, n1303_sel, n920_sel, n546_sel, g158_sel, n1469_sel, n1086_sel, n707_sel, n332_sel, n1252_sel, n869_sel, n495_sel, n1418_sel, n1035_sel, n659_sel, n1201_sel, n807_sel, n447_sel, n1367_sel, n984_sel, n610_sel, n1532_sel, n1150_sel, n762_sel, n396_sel, n1316_sel, n933_sel, n559_sel, n1481_sel, n1099_sel, n4_sel, n345_sel, n1265_sel, n882_sel, n508_sel, n1431_sel, n1048_sel, n672_sel, n1214_sel, n817_sel, n460_sel, n1380_sel, n997_sel, n623_sel, n1545_sel, n1163_sel, n775_sel, n409_sel, n1329_sel, n946_sel, n572_sel, n1494_sel, n1112_sel, n730_sel, n358_sel, n1278_sel, n895_sel, n521_sel, n1444_sel, n1061_sel, n685_sel, n307_sel, n1227_sel, n830_sel, g82_sel, n1393_sel, n1010_sel, n636_sel, n1558_sel, n1176_sel, n785_sel, n422_sel, n1342_sel, n959_sel, n585_sel, n1507_sel, n1125_sel, n740_sel, n371_sel, n1291_sel, n908_sel, n534_sel, g146_sel, n1457_sel, n1074_sel, n698_sel, n320_sel, n1240_sel, n840_sel, n483_sel, g95_sel, n1406_sel, n1023_sel, n647_sel, n1189_sel, n18_sel, n435_sel, n1355_sel, n972_sel, n598_sel, n1520_sel, n1138_sel, n753_sel, n384_sel, n1304_sel, n921_sel, n547_sel, g159_sel, n1470_sel, n1087_sel, n708_sel, n333_sel, n1253_sel, n870_sel, n496_sel, n1419_sel, n1036_sel, n660_sel, n1202_sel, n808_sel, n448_sel, n1368_sel, n985_sel, n611_sel, n1533_sel, n1151_sel, n763_sel, n397_sel, n1317_sel, n934_sel, n560_sel, n1482_sel, n1100_sel, n5_sel, n346_sel, n1266_sel, n883_sel, n509_sel, n1432_sel, n1049_sel, n673_sel, n1215_sel, n818_sel, n461_sel, n1381_sel, n998_sel, n624_sel, n1546_sel, n1164_sel, n776_sel, n410_sel, n1330_sel, n947_sel, n573_sel, n1495_sel, n1113_sel, n731_sel, n359_sel, n1279_sel, n896_sel, n522_sel, n1445_sel, n1062_sel, n686_sel, n308_sel, n1228_sel, n831_sel, n471_sel, g83_sel, n1394_sel, n1011_sel, n637_sel, n1177_sel, n786_sel, n423_sel, n1343_sel, n960_sel, n586_sel, n1508_sel, n1126_sel, n741_sel, n372_sel, n1292_sel, n909_sel, n535_sel, g147_sel, n1458_sel, n1075_sel, n699_sel, n321_sel, n1241_sel, n841_sel, n484_sel, g96_sel, n1407_sel, n1024_sel, n648_sel, n1190_sel, n796_sel, n436_sel, n1356_sel, n973_sel, n599_sel, n1521_sel, n1139_sel, n754_sel, n385_sel, n1305_sel, n922_sel, n548_sel, g160_sel, n1088_sel, n709_sel, n334_sel, n1254_sel, n871_sel, n497_sel, n1420_sel, n1037_sel, n661_sel, n1203_sel, n809_sel, n449_sel, n1369_sel, n986_sel, n612_sel, n1534_sel, n1152_sel, n764_sel, n398_sel, n1318_sel, n935_sel, n561_sel, n1483_sel, n1101_sel, n6_sel, n347_sel, n1267_sel, n884_sel, n510_sel, n1433_sel, n1050_sel, n674_sel, n1216_sel, n819_sel, n462_sel, n1382_sel, n999_sel, n625_sel, n1547_sel, n1165_sel, n13_sel, n411_sel, n1331_sel, n948_sel, n574_sel, n1496_sel, n1114_sel, n732_sel, n360_sel, n1280_sel, n897_sel, n523_sel, n1446_sel, n1063_sel, n687_sel, n309_sel, n1229_sel, n832_sel, n472_sel, g84_sel, n1395_sel, n1012_sel, n1178_sel, n787_sel, n424_sel, n1344_sel, n961_sel, n587_sel, n1509_sel, n1127_sel, n742_sel, n373_sel, n1293_sel, n910_sel, n536_sel, g148_sel, n1459_sel, n1076_sel, n700_sel, n322_sel, n1242_sel, n842_sel, n485_sel, n1408_sel, n1025_sel, n649_sel, n1191_sel, n797_sel, n437_sel, n1357_sel, n974_sel, n600_sel, n1522_sel, n1140_sel, n755_sel, n386_sel, n1306_sel, n923_sel, n549_sel, n1471_sel, n1089_sel, n710_sel, n335_sel, n1255_sel, n872_sel, n498_sel, n1421_sel, n1038_sel, n662_sel, n1204_sel, n810_sel, n450_sel, n1370_sel, n987_sel, n613_sel, n1535_sel, n1153_sel, n765_sel, n399_sel, n1319_sel, n936_sel, n562_sel, n1484_sel, n1102_sel, n720_sel, n348_sel, n1268_sel, n885_sel, n511_sel, n1434_sel, n1051_sel, n675_sel, n1217_sel, n820_sel, n463_sel, n1383_sel, n1000_sel, n626_sel, n1548_sel, n1166_sel, n14_sel, n412_sel, n1332_sel, n949_sel, n575_sel, n1497_sel, n1115_sel, n733_sel, n361_sel, n1281_sel, n898_sel, n524_sel, n1447_sel, n1064_sel, n688_sel, n310_sel, n1230_sel, n833_sel, n473_sel, g85_sel, n1396_sel, n1013_sel, n1179_sel, n425_sel, n788_sel, n1345_sel, n962_sel, n588_sel, n1510_sel, n1128_sel, n374_sel, n743_sel, n1294_sel, n911_sel, n537_sel, g149_sel, n1460_sel, n1077_sel, n323_sel, n701_sel, n1243_sel, n843_sel, n486_sel, n1409_sel, n1026_sel, n650_sel, n1192_sel, n438_sel, n798_sel, n1358_sel, n975_sel, n601_sel, n1523_sel, n1141_sel, n387_sel, n756_sel, n1307_sel, n924_sel, n550_sel, n1472_sel, n1090_sel, n336_sel, n711_sel, n1256_sel, n873_sel, n499_sel, n1422_sel, n1039_sel, n663_sel, n1205_sel, n451_sel, n811_sel, n1371_sel, n988_sel, n614_sel, n1536_sel, n1154_sel, n400_sel, n766_sel, n1320_sel, n937_sel, n563_sel, n1485_sel, n1103_sel, n349_sel, n721_sel, n1269_sel, n886_sel, n512_sel, n1435_sel, n1052_sel, n298_sel, n676_sel, n1218_sel, n821_sel, n464_sel, n1384_sel, n1001_sel, n627_sel, n1549_sel, n1167_sel, n413_sel, n15_sel, n1333_sel, n950_sel, n576_sel, n1498_sel, n1116_sel, n362_sel, n734_sel, n1282_sel, n899_sel, n525_sel, n1448_sel, n1065_sel, n311_sel, n689_sel, n1231_sel, n22_sel, g86_sel, n474_sel, n1397_sel, n1014_sel, n638_sel, n1180_sel, n789_sel, n426_sel, n1346_sel, n963_sel, n589_sel, n1511_sel, n1129_sel, n744_sel, n375_sel, n1295_sel, n912_sel, g150_sel, n538_sel, n1461_sel, n1078_sel, n702_sel, n324_sel, n1244_sel, n844_sel, n487_sel, n1410_sel, n1027_sel, n651_sel, n1193_sel, n799_sel, n439_sel, n1359_sel, n976_sel, n602_sel, n1524_sel, n1142_sel, n757_sel, n388_sel, n1308_sel, n925_sel, n551_sel, n1473_sel, n1091_sel, n712_sel, n337_sel, n1257_sel, n874_sel, n500_sel, n1423_sel, n1040_sel, n664_sel, n1206_sel, n812_sel, n452_sel, n1372_sel, n989_sel, n615_sel, n1537_sel, n1155_sel, n767_sel, n401_sel, n1321_sel, n938_sel, n564_sel, n1486_sel, n1104_sel, n722_sel, n350_sel, n1270_sel, n887_sel, n513_sel, n1436_sel, n1053_sel, n677_sel, n299_sel, n1219_sel, n822_sel, n465_sel, n1385_sel, n1002_sel, n628_sel, n1550_sel, n1168_sel, n777_sel, n414_sel, n1334_sel, n951_sel, n577_sel, n1499_sel, n1117_sel, n735_sel, n363_sel, n1283_sel, n900_sel, n526_sel, n1449_sel, n1066_sel, n690_sel, n312_sel, n1232_sel, n23_sel, n475_sel, g87_sel, n1398_sel, n1015_sel, n639_sel, n1181_sel, n790_sel, n427_sel, n1347_sel, n964_sel, n590_sel, n1512_sel, n1130_sel, n745_sel, n376_sel, n1296_sel, n913_sel, n539_sel, g151_sel, n1462_sel, n1079_sel, n703_sel, n325_sel, n1245_sel, n25_sel, n488_sel, n1411_sel, n1028_sel, n652_sel, n1194_sel, n800_sel, n440_sel, n1360_sel, n977_sel, n603_sel, n1525_sel, n1143_sel, n10_sel, n389_sel, n1309_sel, n926_sel, n552_sel, n1474_sel, n1092_sel, n713_sel, n338_sel, n1258_sel, n875_sel, n501_sel, n1424_sel, n1041_sel, n665_sel, n1207_sel, n813_sel, n453_sel, n1373_sel, n990_sel, n616_sel, n1538_sel, n1156_sel, n768_sel, n402_sel, n1322_sel, n939_sel, n565_sel, n1487_sel, n1105_sel, n723_sel, n351_sel, n1271_sel, n888_sel, n514_sel, n1437_sel, n1054_sel, n678_sel, n300_sel, n1220_sel, n823_sel, n466_sel, n1386_sel, n1003_sel, n629_sel, n1551_sel, n1169_sel, n778_sel, n415_sel, n1335_sel, n952_sel, n578_sel, n1500_sel, n1118_sel, n736_sel, n364_sel, n1284_sel, n901_sel, n527_sel, n1450_sel, n1067_sel, n691_sel, n313_sel, n1233_sel, n24_sel, n476_sel, g88_sel, n1399_sel, n1016_sel, n640_sel, n1182_sel, n791_sel, n428_sel, n1348_sel, n965_sel, n591_sel, n1513_sel, n1131_sel, n746_sel, n377_sel, n1297_sel, n914_sel, n540_sel, g152_sel, n1463_sel, n1080_sel, n704_sel, n326_sel, n1246_sel, n26_sel, n489_sel, n1412_sel, n1029_sel, n653_sel, n1195_sel, n801_sel, n441_sel, n1361_sel, n978_sel, n604_sel, n1526_sel, n1144_sel, n11_sel, n390_sel, n1310_sel, n927_sel, n553_sel, n1475_sel, n1093_sel, n714_sel, n339_sel, n1259_sel, n876_sel, n502_sel, n1425_sel, n1042_sel, n666_sel, n1208_sel, n814_sel, n454_sel, n1374_sel, n991_sel, n617_sel, n1539_sel, n1157_sel, n769_sel, n403_sel, n1323_sel, n940_sel, n566_sel, n1488_sel, n1106_sel, n724_sel, n352_sel, n1272_sel, n889_sel, n515_sel, n1438_sel, n1055_sel, n679_sel, n301_sel, n1221_sel, n824_sel, n467_sel, n1387_sel, n1004_sel, n630_sel, n1552_sel, n1170_sel, n779_sel, n416_sel, n1336_sel, n953_sel, n579_sel, n1501_sel, n1119_sel, n737_sel, n365_sel, n1285_sel, n902_sel, n528_sel, n1451_sel, n1068_sel, n692_sel, n314_sel, n1234_sel, n834_sel, n477_sel, g89_sel, n1400_sel, n1017_sel, n641_sel, n1183_sel, n792_sel, n429_sel;
output g32_po, g33_po, g34_po, g35_po, g36_po, g37_po, g38_po, g39_po, g40_po, g41_po, g42_po, g43_po, g44_po, g45_po, g46_po, g47_po, g48_po, g49_po, g50_po, g51_po, g52_po, g53_po, g54_po, g55_po, g56_po, g57_po, g58_po, g59_po, g60_po, g61_po, g62_po, g63_po, g64_po, g65_po, g66_po, g67_po, g68_po, g69_po, g70_po, g71_po, g72_po, g73_po, g74_po, g75_po, g76_po, g77_po, g78_po, g79_po, g80_po, g81_po, g82_po, g83_po, g84_po, g85_po, g86_po, g87_po, g88_po, g89_po, g90_po, g91_po, g92_po, g93_po, g94_po, g95_po, g96_po, g97_po, g98_po, g99_po, g100_po, g101_po, g102_po, g103_po, g104_po, g105_po, g106_po, g107_po, g108_po, g109_po, g110_po, g111_po, g112_po, g113_po, g114_po, g115_po, g116_po, g117_po, g118_po, g119_po, g120_po, g121_po, g122_po, g123_po, g124_po, g125_po, g126_po, g127_po, g128_po, g129_po, g130_po, g131_po, g132_po, g133_po, g134_po, g135_po, g136_po, g137_po, g138_po, g139_po, g140_po, g141_po, g142_po, g143_po, g144_po, g145_po, g146_po, g147_po, g148_po, g149_po, g150_po, g151_po, g152_po, g153_po, g154_po, g155_po, g156_po, g157_po, g158_po, g159_po, g160_po;
wire g349, g350, g351, g352, g353, g354, g355, g356, g357, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n1, n2, n3, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n4, n5, n6, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n7, n8, n9, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n10, n11, n12, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n13, n14, n15, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n16, n17, n18, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n19, n20, n21, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n22, n23, n24, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n25, n26, n27, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n318_1, n330_1, n339_1, n356_1, n361_1, n365_1, n401_1, n408_1, n415_1, n421_1, n431_1, n438_1, n445_1, n483_1, n495_1, n504_1, n521_1, n526_1, n530_1, n566_1, n573_1, n580_1, n586_1, n596_1, n603_1, n610_1, n689_1, n692_1, n695_1, n698_1, n701_1, n704_1, n727_1, n736_1, n746_1, n755_1, n765_1, n774_1, n784_1, n793_1, n803_1, n812_1, n822_1, n831_1, n838_1, n843_1, n875_1, n883_1, n893_1, n908_1, n915_1, n921_1, n927_1, n936_1, n947_1, n956_1, n964_1, n973_1, n988_1, n992_1, n999_1, n1007_1, n1013_1, n1021_1, n1031_1, n1035_1, n1043_1, n1049_1, n1058_1, n1064_1, n1072_1, n1116_1, n1124_1, n1134_1, n1149_1, n1156_1, n1162_1, n1168_1, n1177_1, n1188_1, n1197_1, n1205_1, n1214_1, n1229_1, n1233_1, n1240_1, n1248_1, n1254_1, n1262_1, n1272_1, n1276_1, n1284_1, n1290_1, n1299_1, n1305_1, n1313_1, n1384_1, n1387_1, n1390_1, n1393_1, n1396_1, n1399_1, n1402_1, n1405_1, n1489_1, n1492_1, n1495_1, n1498_1, n1501_1, n1504_1, n1507_1, n1510_1, g0_mux, g0_xnor, g1_mux, g1_xnor, g2_mux, g2_xnor, g3_mux, g3_xnor, g4_mux, g4_xnor, g5_mux, g5_xnor, g6_mux, g6_xnor, g7_mux, g7_xnor, g8_mux, g8_xnor, g9_mux, g9_xnor, g10_mux, g10_xnor, g11_mux, g11_xnor, g12_mux, g12_xnor, g13_mux, g13_xnor, g14_mux, g14_xnor, g15_mux, g15_xnor, g16_mux, g16_xnor, g17_mux, g17_xnor, g18_mux, g18_xnor, g19_mux, g19_xnor, g20_mux, g20_xnor, g21_mux, g21_xnor, g22_mux, g22_xnor, g23_mux, g23_xnor, g24_mux, g24_xnor, g25_mux, g25_xnor, g26_mux, g26_xnor, g27_mux, g27_xnor, g28_mux, g28_xnor, g29_mux, g29_xnor, g30_mux, g30_xnor, g31_mux, g31_xnor, g349_mux, g349_xnor, g350_mux, g350_xnor, g351_mux, g351_xnor, g352_mux, g352_xnor, g353_mux, g353_xnor, g354_mux, g354_xnor, g355_mux, g355_xnor, g356_mux, g356_xnor, g357_mux, g357_xnor, n28_mux, n28_xnor, n29_mux, n29_xnor, n30_mux, n30_xnor, n31_mux, n31_xnor, n32_mux, n32_xnor, n33_mux, n33_xnor, n34_mux, n34_xnor, n35_mux, n35_xnor, n36_mux, n36_xnor, n37_mux, n37_xnor, n38_mux, n38_xnor, n39_mux, n39_xnor, n40_mux, n40_xnor, n41_mux, n41_xnor, n42_mux, n42_xnor, n43_mux, n43_xnor, n44_mux, n44_xnor, n45_mux, n45_xnor, n46_mux, n46_xnor, n47_mux, n47_xnor, n48_mux, n48_xnor, n49_mux, n49_xnor, n50_mux, n50_xnor, n1349_mux, n1349_xnor, n966_mux, n966_xnor, n592_mux, n592_xnor, n1514_mux, n1514_xnor, n1132_mux, n1132_xnor, n747_mux, n747_xnor, n378_mux, n378_xnor, n1298_mux, n1298_xnor, n915_mux, n915_xnor, n541_mux, n541_xnor, g153_mux, g153_xnor, n1464_mux, n1464_xnor, n1081_mux, n1081_xnor, n705_mux, n705_xnor, n327_mux, n327_xnor, n1247_mux, n1247_xnor, n27_mux, n27_xnor, n490_mux, n490_xnor, n1413_mux, n1413_xnor, n1030_mux, n1030_xnor, n654_mux, n654_xnor, n1196_mux, n1196_xnor, n802_mux, n802_xnor, n442_mux, n442_xnor, n1362_mux, n1362_xnor, n979_mux, n979_xnor, n605_mux, n605_xnor, n1527_mux, n1527_xnor, n1145_mux, n1145_xnor, n12_mux, n12_xnor, n391_mux, n391_xnor, n1311_mux, n1311_xnor, n928_mux, n928_xnor, n554_mux, n554_xnor, n1476_mux, n1476_xnor, n1094_mux, n1094_xnor, n715_mux, n715_xnor, n340_mux, n340_xnor, n1260_mux, n1260_xnor, n877_mux, n877_xnor, n503_mux, n503_xnor, n1426_mux, n1426_xnor, n1043_mux, n1043_xnor, n667_mux, n667_xnor, n1209_mux, n1209_xnor, n19_mux, n19_xnor, n455_mux, n455_xnor, n1375_mux, n1375_xnor, n992_mux, n992_xnor, n618_mux, n618_xnor, n1540_mux, n1540_xnor, n1158_mux, n1158_xnor, n770_mux, n770_xnor, n404_mux, n404_xnor, n1324_mux, n1324_xnor, n941_mux, n941_xnor, n567_mux, n567_xnor, n1489_mux, n1489_xnor, n1107_mux, n1107_xnor, n725_mux, n725_xnor, n353_mux, n353_xnor, n1273_mux, n1273_xnor, n890_mux, n890_xnor, n516_mux, n516_xnor, n1439_mux, n1439_xnor, n1056_mux, n1056_xnor, n680_mux, n680_xnor, n302_mux, n302_xnor, n1222_mux, n1222_xnor, n825_mux, n825_xnor, n468_mux, n468_xnor, n1388_mux, n1388_xnor, n1005_mux, n1005_xnor, n631_mux, n631_xnor, n1553_mux, n1553_xnor, n1171_mux, n1171_xnor, n780_mux, n780_xnor, n417_mux, n417_xnor, n1337_mux, n1337_xnor, n954_mux, n954_xnor, n580_mux, n580_xnor, n1502_mux, n1502_xnor, n1120_mux, n1120_xnor, n738_mux, n738_xnor, n366_mux, n366_xnor, n1286_mux, n1286_xnor, n903_mux, n903_xnor, n529_mux, n529_xnor, n1452_mux, n1452_xnor, n1069_mux, n1069_xnor, n693_mux, n693_xnor, n315_mux, n315_xnor, n1235_mux, n1235_xnor, n835_mux, n835_xnor, n478_mux, n478_xnor, g90_mux, g90_xnor, n1401_mux, n1401_xnor, n1018_mux, n1018_xnor, n642_mux, n642_xnor, n1184_mux, n1184_xnor, n793_mux, n793_xnor, n430_mux, n430_xnor, n1350_mux, n1350_xnor, n967_mux, n967_xnor, n593_mux, n593_xnor, n1515_mux, n1515_xnor, n1133_mux, n1133_xnor, n748_mux, n748_xnor, n379_mux, n379_xnor, n1299_mux, n1299_xnor, n916_mux, n916_xnor, n542_mux, n542_xnor, g154_mux, g154_xnor, n1465_mux, n1465_xnor, n1082_mux, n1082_xnor, n706_mux, n706_xnor, n328_mux, n328_xnor, n1248_mux, n1248_xnor, n845_mux, n845_xnor, n491_mux, n491_xnor, n1414_mux, n1414_xnor, n1031_mux, n1031_xnor, n655_mux, n655_xnor, n1197_mux, n1197_xnor, n803_mux, n803_xnor, n443_mux, n443_xnor, n1363_mux, n1363_xnor, n980_mux, n980_xnor, n606_mux, n606_xnor, n1528_mux, n1528_xnor, n1146_mux, n1146_xnor, n758_mux, n758_xnor, n392_mux, n392_xnor, n1312_mux, n1312_xnor, n929_mux, n929_xnor, n555_mux, n555_xnor, n1477_mux, n1477_xnor, n1095_mux, n1095_xnor, n716_mux, n716_xnor, n341_mux, n341_xnor, n1261_mux, n1261_xnor, n878_mux, n878_xnor, n504_mux, n504_xnor, n1427_mux, n1427_xnor, n1044_mux, n1044_xnor, n668_mux, n668_xnor, n1210_mux, n1210_xnor, n20_mux, n20_xnor, n456_mux, n456_xnor, n1376_mux, n1376_xnor, n993_mux, n993_xnor, n619_mux, n619_xnor, n1541_mux, n1541_xnor, n1159_mux, n1159_xnor, n771_mux, n771_xnor, n405_mux, n405_xnor, n1325_mux, n1325_xnor, n942_mux, n942_xnor, n568_mux, n568_xnor, n1490_mux, n1490_xnor, n1108_mux, n1108_xnor, n726_mux, n726_xnor, n354_mux, n354_xnor, n1274_mux, n1274_xnor, n891_mux, n891_xnor, n517_mux, n517_xnor, n1440_mux, n1440_xnor, n1057_mux, n1057_xnor, n681_mux, n681_xnor, n303_mux, n303_xnor, n1223_mux, n1223_xnor, n826_mux, n826_xnor, n469_mux, n469_xnor, n1389_mux, n1389_xnor, n1006_mux, n1006_xnor, n632_mux, n632_xnor, n1554_mux, n1554_xnor, n1172_mux, n1172_xnor, n781_mux, n781_xnor, n418_mux, n418_xnor, n1338_mux, n1338_xnor, n955_mux, n955_xnor, n581_mux, n581_xnor, n1503_mux, n1503_xnor, n1121_mux, n1121_xnor, n7_mux, n7_xnor, n367_mux, n367_xnor, n1287_mux, n1287_xnor, n904_mux, n904_xnor, n530_mux, n530_xnor, n1453_mux, n1453_xnor, n1070_mux, n1070_xnor, n694_mux, n694_xnor, n316_mux, n316_xnor, n1236_mux, n1236_xnor, n836_mux, n836_xnor, n479_mux, n479_xnor, g91_mux, g91_xnor, n1402_mux, n1402_xnor, n1019_mux, n1019_xnor, n643_mux, n643_xnor, n1185_mux, n1185_xnor, n794_mux, n794_xnor, n431_mux, n431_xnor, n1351_mux, n1351_xnor, n968_mux, n968_xnor, n594_mux, n594_xnor, n1516_mux, n1516_xnor, n1134_mux, n1134_xnor, n749_mux, n749_xnor, n380_mux, n380_xnor, n1300_mux, n1300_xnor, n917_mux, n917_xnor, n543_mux, n543_xnor, g155_mux, g155_xnor, n1466_mux, n1466_xnor, n1083_mux, n1083_xnor, n1_mux, n1_xnor, n329_mux, n329_xnor, n1249_mux, n1249_xnor, n866_mux, n866_xnor, n492_mux, n492_xnor, n1415_mux, n1415_xnor, n1032_mux, n1032_xnor, n656_mux, n656_xnor, n1198_mux, n1198_xnor, n444_mux, n444_xnor, n804_mux, n804_xnor, n1364_mux, n1364_xnor, n981_mux, n981_xnor, n607_mux, n607_xnor, n1529_mux, n1529_xnor, n1147_mux, n1147_xnor, n393_mux, n393_xnor, n759_mux, n759_xnor, n1313_mux, n1313_xnor, n930_mux, n930_xnor, n556_mux, n556_xnor, n1478_mux, n1478_xnor, n1096_mux, n1096_xnor, n717_mux, n717_xnor, n342_mux, n342_xnor, n1262_mux, n1262_xnor, n879_mux, n879_xnor, n505_mux, n505_xnor, n1428_mux, n1428_xnor, n1045_mux, n1045_xnor, n669_mux, n669_xnor, n1211_mux, n1211_xnor, n21_mux, n21_xnor, n457_mux, n457_xnor, n1377_mux, n1377_xnor, n994_mux, n994_xnor, n620_mux, n620_xnor, n1542_mux, n1542_xnor, n1160_mux, n1160_xnor, n406_mux, n406_xnor, n772_mux, n772_xnor, n1326_mux, n1326_xnor, n943_mux, n943_xnor, n569_mux, n569_xnor, n1491_mux, n1491_xnor, n1109_mux, n1109_xnor, n355_mux, n355_xnor, n727_mux, n727_xnor, n1275_mux, n1275_xnor, n892_mux, n892_xnor, n518_mux, n518_xnor, n1441_mux, n1441_xnor, n1058_mux, n1058_xnor, n304_mux, n304_xnor, n682_mux, n682_xnor, n1224_mux, n1224_xnor, n827_mux, n827_xnor, n470_mux, n470_xnor, n1390_mux, n1390_xnor, n1007_mux, n1007_xnor, n633_mux, n633_xnor, n1555_mux, n1555_xnor, n1173_mux, n1173_xnor, n419_mux, n419_xnor, n782_mux, n782_xnor, n1339_mux, n1339_xnor, n956_mux, n956_xnor, n582_mux, n582_xnor, n1504_mux, n1504_xnor, n1122_mux, n1122_xnor, n368_mux, n368_xnor, n8_mux, n8_xnor, n1288_mux, n1288_xnor, n905_mux, n905_xnor, n531_mux, n531_xnor, n1454_mux, n1454_xnor, n1071_mux, n1071_xnor, n317_mux, n317_xnor, n695_mux, n695_xnor, n1237_mux, n1237_xnor, n837_mux, n837_xnor, n480_mux, n480_xnor, g92_mux, g92_xnor, n1403_mux, n1403_xnor, n1020_mux, n1020_xnor, n644_mux, n644_xnor, n1186_mux, n1186_xnor, n432_mux, n432_xnor, n795_mux, n795_xnor, n1352_mux, n1352_xnor, n969_mux, n969_xnor, n595_mux, n595_xnor, n1517_mux, n1517_xnor, n1135_mux, n1135_xnor, n381_mux, n381_xnor, n750_mux, n750_xnor, n1301_mux, n1301_xnor, n918_mux, n918_xnor, g156_mux, g156_xnor, n544_mux, n544_xnor, n1467_mux, n1467_xnor, n1084_mux, n1084_xnor, n330_mux, n330_xnor, n2_mux, n2_xnor, n1250_mux, n1250_xnor, n867_mux, n867_xnor, n493_mux, n493_xnor, n1416_mux, n1416_xnor, n1033_mux, n1033_xnor, n657_mux, n657_xnor, n1199_mux, n1199_xnor, n805_mux, n805_xnor, n445_mux, n445_xnor, n1365_mux, n1365_xnor, n982_mux, n982_xnor, n608_mux, n608_xnor, n1530_mux, n1530_xnor, n1148_mux, n1148_xnor, n760_mux, n760_xnor, n394_mux, n394_xnor, n1314_mux, n1314_xnor, n931_mux, n931_xnor, n557_mux, n557_xnor, n1479_mux, n1479_xnor, n1097_mux, n1097_xnor, n343_mux, n343_xnor, n718_mux, n718_xnor, n1263_mux, n1263_xnor, n880_mux, n880_xnor, n506_mux, n506_xnor, n1429_mux, n1429_xnor, n1046_mux, n1046_xnor, n670_mux, n670_xnor, n1212_mux, n1212_xnor, n815_mux, n815_xnor, n458_mux, n458_xnor, n1378_mux, n1378_xnor, n995_mux, n995_xnor, n621_mux, n621_xnor, n1543_mux, n1543_xnor, n1161_mux, n1161_xnor, n773_mux, n773_xnor, n407_mux, n407_xnor, n1327_mux, n1327_xnor, n944_mux, n944_xnor, n570_mux, n570_xnor, n1492_mux, n1492_xnor, n1110_mux, n1110_xnor, n728_mux, n728_xnor, n356_mux, n356_xnor, n1276_mux, n1276_xnor, n893_mux, n893_xnor, n519_mux, n519_xnor, n1442_mux, n1442_xnor, n1059_mux, n1059_xnor, n683_mux, n683_xnor, n305_mux, n305_xnor, n1225_mux, n1225_xnor, n828_mux, n828_xnor, g80_mux, g80_xnor, n1391_mux, n1391_xnor, n1008_mux, n1008_xnor, n634_mux, n634_xnor, n1556_mux, n1556_xnor, n1174_mux, n1174_xnor, n783_mux, n783_xnor, n420_mux, n420_xnor, n1340_mux, n1340_xnor, n957_mux, n957_xnor, n583_mux, n583_xnor, n1505_mux, n1505_xnor, n1123_mux, n1123_xnor, n9_mux, n9_xnor, n369_mux, n369_xnor, n1289_mux, n1289_xnor, n906_mux, n906_xnor, g144_mux, g144_xnor, n532_mux, n532_xnor, n1455_mux, n1455_xnor, n1072_mux, n1072_xnor, n696_mux, n696_xnor, n318_mux, n318_xnor, n1238_mux, n1238_xnor, n838_mux, n838_xnor, g93_mux, g93_xnor, n481_mux, n481_xnor, n1404_mux, n1404_xnor, n1021_mux, n1021_xnor, n645_mux, n645_xnor, n1187_mux, n1187_xnor, n16_mux, n16_xnor, n433_mux, n433_xnor, n1353_mux, n1353_xnor, n970_mux, n970_xnor, n596_mux, n596_xnor, n1518_mux, n1518_xnor, n1136_mux, n1136_xnor, n751_mux, n751_xnor, n382_mux, n382_xnor, n1302_mux, n1302_xnor, n919_mux, n919_xnor, n545_mux, n545_xnor, g157_mux, g157_xnor, n1468_mux, n1468_xnor, n1085_mux, n1085_xnor, n3_mux, n3_xnor, n331_mux, n331_xnor, n1251_mux, n1251_xnor, n868_mux, n868_xnor, n494_mux, n494_xnor, n1417_mux, n1417_xnor, n1034_mux, n1034_xnor, n658_mux, n658_xnor, n1200_mux, n1200_xnor, n806_mux, n806_xnor, n446_mux, n446_xnor, n1366_mux, n1366_xnor, n983_mux, n983_xnor, n609_mux, n609_xnor, n1531_mux, n1531_xnor, n1149_mux, n1149_xnor, n761_mux, n761_xnor, n395_mux, n395_xnor, n1315_mux, n1315_xnor, n932_mux, n932_xnor, n558_mux, n558_xnor, n1480_mux, n1480_xnor, n1098_mux, n1098_xnor, n719_mux, n719_xnor, n344_mux, n344_xnor, n1264_mux, n1264_xnor, n881_mux, n881_xnor, n507_mux, n507_xnor, n1430_mux, n1430_xnor, n1047_mux, n1047_xnor, n671_mux, n671_xnor, n1213_mux, n1213_xnor, n816_mux, n816_xnor, n459_mux, n459_xnor, n1379_mux, n1379_xnor, n996_mux, n996_xnor, n622_mux, n622_xnor, n1544_mux, n1544_xnor, n1162_mux, n1162_xnor, n774_mux, n774_xnor, n408_mux, n408_xnor, n1328_mux, n1328_xnor, n945_mux, n945_xnor, n571_mux, n571_xnor, n1493_mux, n1493_xnor, n1111_mux, n1111_xnor, n729_mux, n729_xnor, n357_mux, n357_xnor, n1277_mux, n1277_xnor, n894_mux, n894_xnor, n520_mux, n520_xnor, n1443_mux, n1443_xnor, n1060_mux, n1060_xnor, n684_mux, n684_xnor, n306_mux, n306_xnor, n1226_mux, n1226_xnor, n829_mux, n829_xnor, g81_mux, g81_xnor, n1392_mux, n1392_xnor, n1009_mux, n1009_xnor, n635_mux, n635_xnor, n1557_mux, n1557_xnor, n1175_mux, n1175_xnor, n784_mux, n784_xnor, n421_mux, n421_xnor, n1341_mux, n1341_xnor, n958_mux, n958_xnor, n584_mux, n584_xnor, n1506_mux, n1506_xnor, n1124_mux, n1124_xnor, n739_mux, n739_xnor, n370_mux, n370_xnor, n1290_mux, n1290_xnor, n907_mux, n907_xnor, n533_mux, n533_xnor, g145_mux, g145_xnor, n1456_mux, n1456_xnor, n1073_mux, n1073_xnor, n697_mux, n697_xnor, n319_mux, n319_xnor, n1239_mux, n1239_xnor, n839_mux, n839_xnor, n482_mux, n482_xnor, g94_mux, g94_xnor, n1405_mux, n1405_xnor, n1022_mux, n1022_xnor, n646_mux, n646_xnor, n1188_mux, n1188_xnor, n17_mux, n17_xnor, n434_mux, n434_xnor, n1354_mux, n1354_xnor, n971_mux, n971_xnor, n597_mux, n597_xnor, n1519_mux, n1519_xnor, n1137_mux, n1137_xnor, n752_mux, n752_xnor, n383_mux, n383_xnor, n1303_mux, n1303_xnor, n920_mux, n920_xnor, n546_mux, n546_xnor, g158_mux, g158_xnor, n1469_mux, n1469_xnor, n1086_mux, n1086_xnor, n707_mux, n707_xnor, n332_mux, n332_xnor, n1252_mux, n1252_xnor, n869_mux, n869_xnor, n495_mux, n495_xnor, n1418_mux, n1418_xnor, n1035_mux, n1035_xnor, n659_mux, n659_xnor, n1201_mux, n1201_xnor, n807_mux, n807_xnor, n447_mux, n447_xnor, n1367_mux, n1367_xnor, n984_mux, n984_xnor, n610_mux, n610_xnor, n1532_mux, n1532_xnor, n1150_mux, n1150_xnor, n762_mux, n762_xnor, n396_mux, n396_xnor, n1316_mux, n1316_xnor, n933_mux, n933_xnor, n559_mux, n559_xnor, n1481_mux, n1481_xnor, n1099_mux, n1099_xnor, n4_mux, n4_xnor, n345_mux, n345_xnor, n1265_mux, n1265_xnor, n882_mux, n882_xnor, n508_mux, n508_xnor, n1431_mux, n1431_xnor, n1048_mux, n1048_xnor, n672_mux, n672_xnor, n1214_mux, n1214_xnor, n817_mux, n817_xnor, n460_mux, n460_xnor, n1380_mux, n1380_xnor, n997_mux, n997_xnor, n623_mux, n623_xnor, n1545_mux, n1545_xnor, n1163_mux, n1163_xnor, n775_mux, n775_xnor, n409_mux, n409_xnor, n1329_mux, n1329_xnor, n946_mux, n946_xnor, n572_mux, n572_xnor, n1494_mux, n1494_xnor, n1112_mux, n1112_xnor, n730_mux, n730_xnor, n358_mux, n358_xnor, n1278_mux, n1278_xnor, n895_mux, n895_xnor, n521_mux, n521_xnor, n1444_mux, n1444_xnor, n1061_mux, n1061_xnor, n685_mux, n685_xnor, n307_mux, n307_xnor, n1227_mux, n1227_xnor, n830_mux, n830_xnor, g82_mux, g82_xnor, n1393_mux, n1393_xnor, n1010_mux, n1010_xnor, n636_mux, n636_xnor, n1558_mux, n1558_xnor, n1176_mux, n1176_xnor, n785_mux, n785_xnor, n422_mux, n422_xnor, n1342_mux, n1342_xnor, n959_mux, n959_xnor, n585_mux, n585_xnor, n1507_mux, n1507_xnor, n1125_mux, n1125_xnor, n740_mux, n740_xnor, n371_mux, n371_xnor, n1291_mux, n1291_xnor, n908_mux, n908_xnor, n534_mux, n534_xnor, g146_mux, g146_xnor, n1457_mux, n1457_xnor, n1074_mux, n1074_xnor, n698_mux, n698_xnor, n320_mux, n320_xnor, n1240_mux, n1240_xnor, n840_mux, n840_xnor, n483_mux, n483_xnor, g95_mux, g95_xnor, n1406_mux, n1406_xnor, n1023_mux, n1023_xnor, n647_mux, n647_xnor, n1189_mux, n1189_xnor, n18_mux, n18_xnor, n435_mux, n435_xnor, n1355_mux, n1355_xnor, n972_mux, n972_xnor, n598_mux, n598_xnor, n1520_mux, n1520_xnor, n1138_mux, n1138_xnor, n753_mux, n753_xnor, n384_mux, n384_xnor, n1304_mux, n1304_xnor, n921_mux, n921_xnor, n547_mux, n547_xnor, g159_mux, g159_xnor, n1470_mux, n1470_xnor, n1087_mux, n1087_xnor, n708_mux, n708_xnor, n333_mux, n333_xnor, n1253_mux, n1253_xnor, n870_mux, n870_xnor, n496_mux, n496_xnor, n1419_mux, n1419_xnor, n1036_mux, n1036_xnor, n660_mux, n660_xnor, n1202_mux, n1202_xnor, n808_mux, n808_xnor, n448_mux, n448_xnor, n1368_mux, n1368_xnor, n985_mux, n985_xnor, n611_mux, n611_xnor, n1533_mux, n1533_xnor, n1151_mux, n1151_xnor, n763_mux, n763_xnor, n397_mux, n397_xnor, n1317_mux, n1317_xnor, n934_mux, n934_xnor, n560_mux, n560_xnor, n1482_mux, n1482_xnor, n1100_mux, n1100_xnor, n5_mux, n5_xnor, n346_mux, n346_xnor, n1266_mux, n1266_xnor, n883_mux, n883_xnor, n509_mux, n509_xnor, n1432_mux, n1432_xnor, n1049_mux, n1049_xnor, n673_mux, n673_xnor, n1215_mux, n1215_xnor, n818_mux, n818_xnor, n461_mux, n461_xnor, n1381_mux, n1381_xnor, n998_mux, n998_xnor, n624_mux, n624_xnor, n1546_mux, n1546_xnor, n1164_mux, n1164_xnor, n776_mux, n776_xnor, n410_mux, n410_xnor, n1330_mux, n1330_xnor, n947_mux, n947_xnor, n573_mux, n573_xnor, n1495_mux, n1495_xnor, n1113_mux, n1113_xnor, n731_mux, n731_xnor, n359_mux, n359_xnor, n1279_mux, n1279_xnor, n896_mux, n896_xnor, n522_mux, n522_xnor, n1445_mux, n1445_xnor, n1062_mux, n1062_xnor, n686_mux, n686_xnor, n308_mux, n308_xnor, n1228_mux, n1228_xnor, n831_mux, n831_xnor, n471_mux, n471_xnor, g83_mux, g83_xnor, n1394_mux, n1394_xnor, n1011_mux, n1011_xnor, n637_mux, n637_xnor, n1177_mux, n1177_xnor, n786_mux, n786_xnor, n423_mux, n423_xnor, n1343_mux, n1343_xnor, n960_mux, n960_xnor, n586_mux, n586_xnor, n1508_mux, n1508_xnor, n1126_mux, n1126_xnor, n741_mux, n741_xnor, n372_mux, n372_xnor, n1292_mux, n1292_xnor, n909_mux, n909_xnor, n535_mux, n535_xnor, g147_mux, g147_xnor, n1458_mux, n1458_xnor, n1075_mux, n1075_xnor, n699_mux, n699_xnor, n321_mux, n321_xnor, n1241_mux, n1241_xnor, n841_mux, n841_xnor, n484_mux, n484_xnor, g96_mux, g96_xnor, n1407_mux, n1407_xnor, n1024_mux, n1024_xnor, n648_mux, n648_xnor, n1190_mux, n1190_xnor, n796_mux, n796_xnor, n436_mux, n436_xnor, n1356_mux, n1356_xnor, n973_mux, n973_xnor, n599_mux, n599_xnor, n1521_mux, n1521_xnor, n1139_mux, n1139_xnor, n754_mux, n754_xnor, n385_mux, n385_xnor, n1305_mux, n1305_xnor, n922_mux, n922_xnor, n548_mux, n548_xnor, g160_mux, g160_xnor, n1088_mux, n1088_xnor, n709_mux, n709_xnor, n334_mux, n334_xnor, n1254_mux, n1254_xnor, n871_mux, n871_xnor, n497_mux, n497_xnor, n1420_mux, n1420_xnor, n1037_mux, n1037_xnor, n661_mux, n661_xnor, n1203_mux, n1203_xnor, n809_mux, n809_xnor, n449_mux, n449_xnor, n1369_mux, n1369_xnor, n986_mux, n986_xnor, n612_mux, n612_xnor, n1534_mux, n1534_xnor, n1152_mux, n1152_xnor, n764_mux, n764_xnor, n398_mux, n398_xnor, n1318_mux, n1318_xnor, n935_mux, n935_xnor, n561_mux, n561_xnor, n1483_mux, n1483_xnor, n1101_mux, n1101_xnor, n6_mux, n6_xnor, n347_mux, n347_xnor, n1267_mux, n1267_xnor, n884_mux, n884_xnor, n510_mux, n510_xnor, n1433_mux, n1433_xnor, n1050_mux, n1050_xnor, n674_mux, n674_xnor, n1216_mux, n1216_xnor, n819_mux, n819_xnor, n462_mux, n462_xnor, n1382_mux, n1382_xnor, n999_mux, n999_xnor, n625_mux, n625_xnor, n1547_mux, n1547_xnor, n1165_mux, n1165_xnor, n13_mux, n13_xnor, n411_mux, n411_xnor, n1331_mux, n1331_xnor, n948_mux, n948_xnor, n574_mux, n574_xnor, n1496_mux, n1496_xnor, n1114_mux, n1114_xnor, n732_mux, n732_xnor, n360_mux, n360_xnor, n1280_mux, n1280_xnor, n897_mux, n897_xnor, n523_mux, n523_xnor, n1446_mux, n1446_xnor, n1063_mux, n1063_xnor, n687_mux, n687_xnor, n309_mux, n309_xnor, n1229_mux, n1229_xnor, n832_mux, n832_xnor, n472_mux, n472_xnor, g84_mux, g84_xnor, n1395_mux, n1395_xnor, n1012_mux, n1012_xnor, n1178_mux, n1178_xnor, n787_mux, n787_xnor, n424_mux, n424_xnor, n1344_mux, n1344_xnor, n961_mux, n961_xnor, n587_mux, n587_xnor, n1509_mux, n1509_xnor, n1127_mux, n1127_xnor, n742_mux, n742_xnor, n373_mux, n373_xnor, n1293_mux, n1293_xnor, n910_mux, n910_xnor, n536_mux, n536_xnor, g148_mux, g148_xnor, n1459_mux, n1459_xnor, n1076_mux, n1076_xnor, n700_mux, n700_xnor, n322_mux, n322_xnor, n1242_mux, n1242_xnor, n842_mux, n842_xnor, n485_mux, n485_xnor, n1408_mux, n1408_xnor, n1025_mux, n1025_xnor, n649_mux, n649_xnor, n1191_mux, n1191_xnor, n797_mux, n797_xnor, n437_mux, n437_xnor, n1357_mux, n1357_xnor, n974_mux, n974_xnor, n600_mux, n600_xnor, n1522_mux, n1522_xnor, n1140_mux, n1140_xnor, n755_mux, n755_xnor, n386_mux, n386_xnor, n1306_mux, n1306_xnor, n923_mux, n923_xnor, n549_mux, n549_xnor, n1471_mux, n1471_xnor, n1089_mux, n1089_xnor, n710_mux, n710_xnor, n335_mux, n335_xnor, n1255_mux, n1255_xnor, n872_mux, n872_xnor, n498_mux, n498_xnor, n1421_mux, n1421_xnor, n1038_mux, n1038_xnor, n662_mux, n662_xnor, n1204_mux, n1204_xnor, n810_mux, n810_xnor, n450_mux, n450_xnor, n1370_mux, n1370_xnor, n987_mux, n987_xnor, n613_mux, n613_xnor, n1535_mux, n1535_xnor, n1153_mux, n1153_xnor, n765_mux, n765_xnor, n399_mux, n399_xnor, n1319_mux, n1319_xnor, n936_mux, n936_xnor, n562_mux, n562_xnor, n1484_mux, n1484_xnor, n1102_mux, n1102_xnor, n720_mux, n720_xnor, n348_mux, n348_xnor, n1268_mux, n1268_xnor, n885_mux, n885_xnor, n511_mux, n511_xnor, n1434_mux, n1434_xnor, n1051_mux, n1051_xnor, n675_mux, n675_xnor, n1217_mux, n1217_xnor, n820_mux, n820_xnor, n463_mux, n463_xnor, n1383_mux, n1383_xnor, n1000_mux, n1000_xnor, n626_mux, n626_xnor, n1548_mux, n1548_xnor, n1166_mux, n1166_xnor, n14_mux, n14_xnor, n412_mux, n412_xnor, n1332_mux, n1332_xnor, n949_mux, n949_xnor, n575_mux, n575_xnor, n1497_mux, n1497_xnor, n1115_mux, n1115_xnor, n733_mux, n733_xnor, n361_mux, n361_xnor, n1281_mux, n1281_xnor, n898_mux, n898_xnor, n524_mux, n524_xnor, n1447_mux, n1447_xnor, n1064_mux, n1064_xnor, n688_mux, n688_xnor, n310_mux, n310_xnor, n1230_mux, n1230_xnor, n833_mux, n833_xnor, n473_mux, n473_xnor, g85_mux, g85_xnor, n1396_mux, n1396_xnor, n1013_mux, n1013_xnor, n1179_mux, n1179_xnor, n425_mux, n425_xnor, n788_mux, n788_xnor, n1345_mux, n1345_xnor, n962_mux, n962_xnor, n588_mux, n588_xnor, n1510_mux, n1510_xnor, n1128_mux, n1128_xnor, n374_mux, n374_xnor, n743_mux, n743_xnor, n1294_mux, n1294_xnor, n911_mux, n911_xnor, n537_mux, n537_xnor, g149_mux, g149_xnor, n1460_mux, n1460_xnor, n1077_mux, n1077_xnor, n323_mux, n323_xnor, n701_mux, n701_xnor, n1243_mux, n1243_xnor, n843_mux, n843_xnor, n486_mux, n486_xnor, n1409_mux, n1409_xnor, n1026_mux, n1026_xnor, n650_mux, n650_xnor, n1192_mux, n1192_xnor, n438_mux, n438_xnor, n798_mux, n798_xnor, n1358_mux, n1358_xnor, n975_mux, n975_xnor, n601_mux, n601_xnor, n1523_mux, n1523_xnor, n1141_mux, n1141_xnor, n387_mux, n387_xnor, n756_mux, n756_xnor, n1307_mux, n1307_xnor, n924_mux, n924_xnor, n550_mux, n550_xnor, n1472_mux, n1472_xnor, n1090_mux, n1090_xnor, n336_mux, n336_xnor, n711_mux, n711_xnor, n1256_mux, n1256_xnor, n873_mux, n873_xnor, n499_mux, n499_xnor, n1422_mux, n1422_xnor, n1039_mux, n1039_xnor, n663_mux, n663_xnor, n1205_mux, n1205_xnor, n451_mux, n451_xnor, n811_mux, n811_xnor, n1371_mux, n1371_xnor, n988_mux, n988_xnor, n614_mux, n614_xnor, n1536_mux, n1536_xnor, n1154_mux, n1154_xnor, n400_mux, n400_xnor, n766_mux, n766_xnor, n1320_mux, n1320_xnor, n937_mux, n937_xnor, n563_mux, n563_xnor, n1485_mux, n1485_xnor, n1103_mux, n1103_xnor, n349_mux, n349_xnor, n721_mux, n721_xnor, n1269_mux, n1269_xnor, n886_mux, n886_xnor, n512_mux, n512_xnor, n1435_mux, n1435_xnor, n1052_mux, n1052_xnor, n298_mux, n298_xnor, n676_mux, n676_xnor, n1218_mux, n1218_xnor, n821_mux, n821_xnor, n464_mux, n464_xnor, n1384_mux, n1384_xnor, n1001_mux, n1001_xnor, n627_mux, n627_xnor, n1549_mux, n1549_xnor, n1167_mux, n1167_xnor, n413_mux, n413_xnor, n15_mux, n15_xnor, n1333_mux, n1333_xnor, n950_mux, n950_xnor, n576_mux, n576_xnor, n1498_mux, n1498_xnor, n1116_mux, n1116_xnor, n362_mux, n362_xnor, n734_mux, n734_xnor, n1282_mux, n1282_xnor, n899_mux, n899_xnor, n525_mux, n525_xnor, n1448_mux, n1448_xnor, n1065_mux, n1065_xnor, n311_mux, n311_xnor, n689_mux, n689_xnor, n1231_mux, n1231_xnor, n22_mux, n22_xnor, g86_mux, g86_xnor, n474_mux, n474_xnor, n1397_mux, n1397_xnor, n1014_mux, n1014_xnor, n638_mux, n638_xnor, n1180_mux, n1180_xnor, n789_mux, n789_xnor, n426_mux, n426_xnor, n1346_mux, n1346_xnor, n963_mux, n963_xnor, n589_mux, n589_xnor, n1511_mux, n1511_xnor, n1129_mux, n1129_xnor, n744_mux, n744_xnor, n375_mux, n375_xnor, n1295_mux, n1295_xnor, n912_mux, n912_xnor, g150_mux, g150_xnor, n538_mux, n538_xnor, n1461_mux, n1461_xnor, n1078_mux, n1078_xnor, n702_mux, n702_xnor, n324_mux, n324_xnor, n1244_mux, n1244_xnor, n844_mux, n844_xnor, n487_mux, n487_xnor, n1410_mux, n1410_xnor, n1027_mux, n1027_xnor, n651_mux, n651_xnor, n1193_mux, n1193_xnor, n799_mux, n799_xnor, n439_mux, n439_xnor, n1359_mux, n1359_xnor, n976_mux, n976_xnor, n602_mux, n602_xnor, n1524_mux, n1524_xnor, n1142_mux, n1142_xnor, n757_mux, n757_xnor, n388_mux, n388_xnor, n1308_mux, n1308_xnor, n925_mux, n925_xnor, n551_mux, n551_xnor, n1473_mux, n1473_xnor, n1091_mux, n1091_xnor, n712_mux, n712_xnor, n337_mux, n337_xnor, n1257_mux, n1257_xnor, n874_mux, n874_xnor, n500_mux, n500_xnor, n1423_mux, n1423_xnor, n1040_mux, n1040_xnor, n664_mux, n664_xnor, n1206_mux, n1206_xnor, n812_mux, n812_xnor, n452_mux, n452_xnor, n1372_mux, n1372_xnor, n989_mux, n989_xnor, n615_mux, n615_xnor, n1537_mux, n1537_xnor, n1155_mux, n1155_xnor, n767_mux, n767_xnor, n401_mux, n401_xnor, n1321_mux, n1321_xnor, n938_mux, n938_xnor, n564_mux, n564_xnor, n1486_mux, n1486_xnor, n1104_mux, n1104_xnor, n722_mux, n722_xnor, n350_mux, n350_xnor, n1270_mux, n1270_xnor, n887_mux, n887_xnor, n513_mux, n513_xnor, n1436_mux, n1436_xnor, n1053_mux, n1053_xnor, n677_mux, n677_xnor, n299_mux, n299_xnor, n1219_mux, n1219_xnor, n822_mux, n822_xnor, n465_mux, n465_xnor, n1385_mux, n1385_xnor, n1002_mux, n1002_xnor, n628_mux, n628_xnor, n1550_mux, n1550_xnor, n1168_mux, n1168_xnor, n777_mux, n777_xnor, n414_mux, n414_xnor, n1334_mux, n1334_xnor, n951_mux, n951_xnor, n577_mux, n577_xnor, n1499_mux, n1499_xnor, n1117_mux, n1117_xnor, n735_mux, n735_xnor, n363_mux, n363_xnor, n1283_mux, n1283_xnor, n900_mux, n900_xnor, n526_mux, n526_xnor, n1449_mux, n1449_xnor, n1066_mux, n1066_xnor, n690_mux, n690_xnor, n312_mux, n312_xnor, n1232_mux, n1232_xnor, n23_mux, n23_xnor, n475_mux, n475_xnor, g87_mux, g87_xnor, n1398_mux, n1398_xnor, n1015_mux, n1015_xnor, n639_mux, n639_xnor, n1181_mux, n1181_xnor, n790_mux, n790_xnor, n427_mux, n427_xnor, n1347_mux, n1347_xnor, n964_mux, n964_xnor, n590_mux, n590_xnor, n1512_mux, n1512_xnor, n1130_mux, n1130_xnor, n745_mux, n745_xnor, n376_mux, n376_xnor, n1296_mux, n1296_xnor, n913_mux, n913_xnor, n539_mux, n539_xnor, g151_mux, g151_xnor, n1462_mux, n1462_xnor, n1079_mux, n1079_xnor, n703_mux, n703_xnor, n325_mux, n325_xnor, n1245_mux, n1245_xnor, n25_mux, n25_xnor, n488_mux, n488_xnor, n1411_mux, n1411_xnor, n1028_mux, n1028_xnor, n652_mux, n652_xnor, n1194_mux, n1194_xnor, n800_mux, n800_xnor, n440_mux, n440_xnor, n1360_mux, n1360_xnor, n977_mux, n977_xnor, n603_mux, n603_xnor, n1525_mux, n1525_xnor, n1143_mux, n1143_xnor, n10_mux, n10_xnor, n389_mux, n389_xnor, n1309_mux, n1309_xnor, n926_mux, n926_xnor, n552_mux, n552_xnor, n1474_mux, n1474_xnor, n1092_mux, n1092_xnor, n713_mux, n713_xnor, n338_mux, n338_xnor, n1258_mux, n1258_xnor, n875_mux, n875_xnor, n501_mux, n501_xnor, n1424_mux, n1424_xnor, n1041_mux, n1041_xnor, n665_mux, n665_xnor, n1207_mux, n1207_xnor, n813_mux, n813_xnor, n453_mux, n453_xnor, n1373_mux, n1373_xnor, n990_mux, n990_xnor, n616_mux, n616_xnor, n1538_mux, n1538_xnor, n1156_mux, n1156_xnor, n768_mux, n768_xnor, n402_mux, n402_xnor, n1322_mux, n1322_xnor, n939_mux, n939_xnor, n565_mux, n565_xnor, n1487_mux, n1487_xnor, n1105_mux, n1105_xnor, n723_mux, n723_xnor, n351_mux, n351_xnor, n1271_mux, n1271_xnor, n888_mux, n888_xnor, n514_mux, n514_xnor, n1437_mux, n1437_xnor, n1054_mux, n1054_xnor, n678_mux, n678_xnor, n300_mux, n300_xnor, n1220_mux, n1220_xnor, n823_mux, n823_xnor, n466_mux, n466_xnor, n1386_mux, n1386_xnor, n1003_mux, n1003_xnor, n629_mux, n629_xnor, n1551_mux, n1551_xnor, n1169_mux, n1169_xnor, n778_mux, n778_xnor, n415_mux, n415_xnor, n1335_mux, n1335_xnor, n952_mux, n952_xnor, n578_mux, n578_xnor, n1500_mux, n1500_xnor, n1118_mux, n1118_xnor, n736_mux, n736_xnor, n364_mux, n364_xnor, n1284_mux, n1284_xnor, n901_mux, n901_xnor, n527_mux, n527_xnor, n1450_mux, n1450_xnor, n1067_mux, n1067_xnor, n691_mux, n691_xnor, n313_mux, n313_xnor, n1233_mux, n1233_xnor, n24_mux, n24_xnor, n476_mux, n476_xnor, g88_mux, g88_xnor, n1399_mux, n1399_xnor, n1016_mux, n1016_xnor, n640_mux, n640_xnor, n1182_mux, n1182_xnor, n791_mux, n791_xnor, n428_mux, n428_xnor, n1348_mux, n1348_xnor, n965_mux, n965_xnor, n591_mux, n591_xnor, n1513_mux, n1513_xnor, n1131_mux, n1131_xnor, n746_mux, n746_xnor, n377_mux, n377_xnor, n1297_mux, n1297_xnor, n914_mux, n914_xnor, n540_mux, n540_xnor, g152_mux, g152_xnor, n1463_mux, n1463_xnor, n1080_mux, n1080_xnor, n704_mux, n704_xnor, n326_mux, n326_xnor, n1246_mux, n1246_xnor, n26_mux, n26_xnor, n489_mux, n489_xnor, n1412_mux, n1412_xnor, n1029_mux, n1029_xnor, n653_mux, n653_xnor, n1195_mux, n1195_xnor, n801_mux, n801_xnor, n441_mux, n441_xnor, n1361_mux, n1361_xnor, n978_mux, n978_xnor, n604_mux, n604_xnor, n1526_mux, n1526_xnor, n1144_mux, n1144_xnor, n11_mux, n11_xnor, n390_mux, n390_xnor, n1310_mux, n1310_xnor, n927_mux, n927_xnor, n553_mux, n553_xnor, n1475_mux, n1475_xnor, n1093_mux, n1093_xnor, n714_mux, n714_xnor, n339_mux, n339_xnor, n1259_mux, n1259_xnor, n876_mux, n876_xnor, n502_mux, n502_xnor, n1425_mux, n1425_xnor, n1042_mux, n1042_xnor, n666_mux, n666_xnor, n1208_mux, n1208_xnor, n814_mux, n814_xnor, n454_mux, n454_xnor, n1374_mux, n1374_xnor, n991_mux, n991_xnor, n617_mux, n617_xnor, n1539_mux, n1539_xnor, n1157_mux, n1157_xnor, n769_mux, n769_xnor, n403_mux, n403_xnor, n1323_mux, n1323_xnor, n940_mux, n940_xnor, n566_mux, n566_xnor, n1488_mux, n1488_xnor, n1106_mux, n1106_xnor, n724_mux, n724_xnor, n352_mux, n352_xnor, n1272_mux, n1272_xnor, n889_mux, n889_xnor, n515_mux, n515_xnor, n1438_mux, n1438_xnor, n1055_mux, n1055_xnor, n679_mux, n679_xnor, n301_mux, n301_xnor, n1221_mux, n1221_xnor, n824_mux, n824_xnor, n467_mux, n467_xnor, n1387_mux, n1387_xnor, n1004_mux, n1004_xnor, n630_mux, n630_xnor, n1552_mux, n1552_xnor, n1170_mux, n1170_xnor, n779_mux, n779_xnor, n416_mux, n416_xnor, n1336_mux, n1336_xnor, n953_mux, n953_xnor, n579_mux, n579_xnor, n1501_mux, n1501_xnor, n1119_mux, n1119_xnor, n737_mux, n737_xnor, n365_mux, n365_xnor, n1285_mux, n1285_xnor, n902_mux, n902_xnor, n528_mux, n528_xnor, n1451_mux, n1451_xnor, n1068_mux, n1068_xnor, n692_mux, n692_xnor, n314_mux, n314_xnor, n1234_mux, n1234_xnor, n834_mux, n834_xnor, n477_mux, n477_xnor, g89_mux, g89_xnor, n1400_mux, n1400_xnor, n1017_mux, n1017_xnor, n641_mux, n641_xnor, n1183_mux, n1183_xnor, n792_mux, n792_xnor, n429_mux, n429_xnor;
wire t_0, t_1;
buf(n51, 1'b0);
buf(g32, n51);
buf(n52, 1'b0);
buf(g33, n52);
buf(n53, 1'b0);
buf(g34, n53);
buf(n54, 1'b0);
buf(g35, n54);
buf(n55, 1'b0);
buf(g36, n55);
buf(n56, 1'b0);
buf(g37, n56);
buf(n57, 1'b0);
buf(g38, n57);
buf(n58, 1'b0);
buf(g39, n58);
buf(n59, 1'b0);
buf(g40, n59);
buf(n60, 1'b0);
buf(g41, n60);
buf(n61, 1'b0);
buf(g42, n61);
buf(n62, 1'b0);
buf(g43, n62);
buf(n63, 1'b0);
buf(g44, n63);
buf(n64, 1'b0);
buf(g45, n64);
buf(n65, 1'b0);
buf(g46, n65);
buf(n66, 1'b0);
buf(g47, n66);
buf(n67, 1'b0);
buf(g48, n67);
buf(n68, 1'b0);
buf(g49, n68);
buf(n69, 1'b0);
buf(g50, n69);
buf(n70, 1'b0);
buf(g51, n70);
buf(n71, 1'b0);
buf(g52, n71);
buf(n72, 1'b0);
buf(g53, n72);
buf(n73, 1'b0);
buf(g54, n73);
buf(n74, 1'b0);
buf(g55, n74);
buf(n75, 1'b0);
buf(g56, n75);
buf(n76, 1'b0);
buf(g57, n76);
buf(n77, 1'b0);
buf(g58, n77);
buf(n78, 1'b0);
buf(g59, n78);
buf(n79, 1'b0);
buf(g60, n79);
buf(n80, 1'b0);
buf(g61, n80);
buf(n81, 1'b0);
buf(g62, n81);
buf(n82, 1'b0);
buf(g63, n82);
buf(n83, 1'b0);
buf(g64, n83);
buf(n84, 1'b0);
buf(g65, n84);
buf(n85, 1'b0);
buf(g66, n85);
buf(n86, 1'b0);
buf(g67, n86);
buf(n87, 1'b0);
buf(g68, n87);
buf(n88, 1'b0);
buf(g69, n88);
buf(n89, 1'b0);
buf(g70, n89);
buf(n90, 1'b0);
buf(g71, n90);
buf(n91, 1'b0);
buf(g72, n91);
buf(n92, 1'b0);
buf(g73, n92);
buf(n93, 1'b0);
buf(g74, n93);
buf(n94, 1'b0);
buf(g75, n94);
buf(n95, 1'b0);
buf(g76, n95);
buf(n96, 1'b0);
buf(g77, n96);
buf(n97, 1'b0);
buf(g78, n97);
buf(n98, 1'b0);
buf(g79, n98);
buf(g349, g0_mux);
buf(n384, g349_mux);
buf(n35, g16_mux);
buf(n380, n35_mux);
and (n1107, n384_mux, n380_mux);
buf(g352, g3_mux);
buf(n325, g352_mux);
not(n1108, n325_mux);
not(n381, n380_mux);
and (n1109, n381_mux, n325_mux);
nor (n1110, n1108_mux, n1109_mux);
buf(g351, g2_mux);
buf(n334, g351_mux);
buf(n36, g17_mux);
buf(n307, n36_mux);
and (n1111, n334_mux, n307_mux);
and (n1112, n1110_mux, n1111_mux);
buf(g350, g1_mux);
buf(n350, g350_mux);
buf(n37, g18_mux);
buf(n310, n37_mux);
and (n1113, n350_mux, n310_mux);
and (n1114, n1111_mux, n1113_mux);
and (n1115, n1110_mux, n1113_mux);
or (n1116_1, n1114_mux, n1115_mux);
or (n1116, n1112_mux, n1116_1);
not(n1117, n334_mux);
and (n1118, n381_mux, n334_mux);
nor (n1119, n1117_mux, n1118_mux);
and (n1120, n1116_mux, n1119_mux);
and (n1121, n350_mux, n307_mux);
and (n1122, n1119_mux, n1121_mux);
and (n1123, n1116_mux, n1121_mux);
or (n1124_1, n1122_mux, n1123_mux);
or (n1124, n1120_mux, n1124_1);
not(n1125, n350_mux);
and (n1126, n381_mux, n350_mux);
nor (n1127, n1125_mux, n1126_mux);
and (n1128, n1124_mux, n1127_mux);
not(n385, n384_mux);
and (n1129, n385_mux, n307_mux);
not(n1130, n307_mux);
nor (n1131, n1129_mux, n1130_mux);
and (n1132, n1127_mux, n1131_mux);
and (n1133, n1124_mux, n1131_mux);
or (n1134_1, n1132_mux, n1133_mux);
or (n1134, n1128_mux, n1134_1);
and (n1135, n1107_mux, n1134_mux);
xor (n1136, n1107_mux, n1134_mux);
xor (n1137, n1124_mux, n1127_mux);
xor (n1138, n1137_mux, n1131_mux);
buf(g353, g4_mux);
buf(n321, g353_mux);
not(n1139, n321_mux);
and (n1140, n381_mux, n321_mux);
nor (n1141, n1139_mux, n1140_mux);
and (n1142, n325_mux, n307_mux);
and (n1143, n1141_mux, n1142_mux);
buf(n39, g20_mux);
buf(n344, n39_mux);
and (n1144, n385_mux, n344_mux);
not(n1145, n344_mux);
nor (n1146, n1144_mux, n1145_mux);
and (n1147, n1142_mux, n1146_mux);
and (n1148, n1141_mux, n1146_mux);
or (n1149_1, n1147_mux, n1148_mux);
or (n1149, n1143_mux, n1149_1);
and (n1150, n325_mux, n310_mux);
buf(n38, g19_mux);
buf(n314, n38_mux);
and (n1151, n334_mux, n314_mux);
and (n1152, n1150_mux, n1151_mux);
and (n1153, n350_mux, n344_mux);
and (n1154, n1151_mux, n1153_mux);
and (n1155, n1150_mux, n1153_mux);
or (n1156_1, n1154_mux, n1155_mux);
or (n1156, n1152_mux, n1156_1);
and (n1157, n334_mux, n310_mux);
and (n1158, n1156_mux, n1157_mux);
and (n1159, n350_mux, n314_mux);
and (n1160, n1157_mux, n1159_mux);
and (n1161, n1156_mux, n1159_mux);
or (n1162_1, n1160_mux, n1161_mux);
or (n1162, n1158_mux, n1162_1);
and (n1163, n1149_mux, n1162_mux);
xor (n1164, n1110_mux, n1111_mux);
xor (n1165, n1164_mux, n1113_mux);
and (n1166, n1162_mux, n1165_mux);
and (n1167, n1149_mux, n1165_mux);
or (n1168_1, n1166_mux, n1167_mux);
or (n1168, n1163_mux, n1168_1);
and (n1169, n385_mux, n310_mux);
not(n1170, n310_mux);
nor (n1171, n1169_mux, n1170_mux);
and (n1172, n1168_mux, n1171_mux);
xor (n1173, n1116_mux, n1119_mux);
xor (n1174, n1173_mux, n1121_mux);
and (n1175, n1171_mux, n1174_mux);
and (n1176, n1168_mux, n1174_mux);
or (n1177_1, n1175_mux, n1176_mux);
or (n1177, n1172_mux, n1177_1);
and (n1178, n1138_mux, n1177_mux);
xor (n1179, n1138_mux, n1177_mux);
xor (n1180, n1168_mux, n1171_mux);
xor (n1181, n1180_mux, n1174_mux);
and (n1182, n325_mux, n314_mux);
and (n1183, n334_mux, n344_mux);
and (n1184, n1182_mux, n1183_mux);
buf(n40, g21_mux);
buf(n319, n40_mux);
and (n1185, n350_mux, n319_mux);
and (n1186, n1183_mux, n1185_mux);
and (n1187, n1182_mux, n1185_mux);
or (n1188_1, n1186_mux, n1187_mux);
or (n1188, n1184_mux, n1188_1);
buf(g354, g5_mux);
buf(n313, g354_mux);
and (n1189, n313_mux, n307_mux);
and (n1190, n321_mux, n310_mux);
and (n1191, n1189_mux, n1190_mux);
and (n1192, n1188_mux, n1191_mux);
xor (n1193, n1150_mux, n1151_mux);
xor (n1194, n1193_mux, n1153_mux);
and (n1195, n1191_mux, n1194_mux);
and (n1196, n1188_mux, n1194_mux);
or (n1197_1, n1195_mux, n1196_mux);
or (n1197, n1192_mux, n1197_1);
xor (n1198, n1141_mux, n1142_mux);
xor (n1199, n1198_mux, n1146_mux);
and (n1200, n1197_mux, n1199_mux);
xor (n1201, n1156_mux, n1157_mux);
xor (n1202, n1201_mux, n1159_mux);
and (n1203, n1199_mux, n1202_mux);
and (n1204, n1197_mux, n1202_mux);
or (n1205_1, n1203_mux, n1204_mux);
or (n1205, n1200_mux, n1205_1);
and (n1206, n385_mux, n314_mux);
not(n1207, n314_mux);
nor (n1208, n1206_mux, n1207_mux);
and (n1209, n1205_mux, n1208_mux);
xor (n1210, n1149_mux, n1162_mux);
xor (n1211, n1210_mux, n1165_mux);
and (n1212, n1208_mux, n1211_mux);
and (n1213, n1205_mux, n1211_mux);
or (n1214_1, n1212_mux, n1213_mux);
or (n1214, n1209_mux, n1214_1);
and (n1215, n1181_mux, n1214_mux);
xor (n1216, n1181_mux, n1214_mux);
xor (n1217, n1205_mux, n1208_mux);
xor (n1218, n1217_mux, n1211_mux);
not(n1219, n313_mux);
and (n1220, n381_mux, n313_mux);
nor (n1221, n1219_mux, n1220_mux);
and (n1222, n321_mux, n307_mux);
and (n1223, n1221_mux, n1222_mux);
and (n1224, n385_mux, n319_mux);
not(n1225, n319_mux);
nor (n1226, n1224_mux, n1225_mux);
and (n1227, n1222_mux, n1226_mux);
and (n1228, n1221_mux, n1226_mux);
or (n1229_1, n1227_mux, n1228_mux);
or (n1229, n1223_mux, n1229_1);
and (n372, n325_mux, n344_mux);
and (n373, n334_mux, n319_mux);
and (n1230, n372_mux, n373_mux);
buf(n41, g22_mux);
buf(n322, n41_mux);
and (n375, n350_mux, n322_mux);
and (n1231, n373_mux, n375_mux);
and (n1232, n372_mux, n375_mux);
or (n1233_1, n1231_mux, n1232_mux);
or (n1233, n1230_mux, n1233_1);
xor (n1234, n1182_mux, n1183_mux);
xor (n1235, n1234_mux, n1185_mux);
and (n1236, n1233_mux, n1235_mux);
xor (n1237, n1189_mux, n1190_mux);
and (n1238, n1235_mux, n1237_mux);
and (n1239, n1233_mux, n1237_mux);
or (n1240_1, n1238_mux, n1239_mux);
or (n1240, n1236_mux, n1240_1);
xor (n1241, n1221_mux, n1222_mux);
xor (n1242, n1241_mux, n1226_mux);
and (n1243, n1240_mux, n1242_mux);
xor (n1244, n1188_mux, n1191_mux);
xor (n1245, n1244_mux, n1194_mux);
and (n1246, n1242_mux, n1245_mux);
and (n1247, n1240_mux, n1245_mux);
or (n1248_1, n1246_mux, n1247_mux);
or (n1248, n1243_mux, n1248_1);
and (n1249, n1229_mux, n1248_mux);
xor (n1250, n1197_mux, n1199_mux);
xor (n1251, n1250_mux, n1202_mux);
and (n1252, n1248_mux, n1251_mux);
and (n1253, n1229_mux, n1251_mux);
or (n1254_1, n1252_mux, n1253_mux);
or (n1254, n1249_mux, n1254_1);
and (n1255, n1218_mux, n1254_mux);
xor (n1256, n1218_mux, n1254_mux);
xor (n1257, n1229_mux, n1248_mux);
xor (n1258, n1257_mux, n1251_mux);
buf(g355, g6_mux);
buf(n309, g355_mux);
and (n366, n309_mux, n307_mux);
and (n367, n313_mux, n310_mux);
and (n1259, n366_mux, n367_mux);
and (n369, n321_mux, n314_mux);
and (n1260, n367_mux, n369_mux);
and (n1261, n366_mux, n369_mux);
or (n1262_1, n1260_mux, n1261_mux);
or (n1262, n1259_mux, n1262_1);
not(n1263, n309_mux);
and (n1264, n381_mux, n309_mux);
nor (n1265, n1263_mux, n1264_mux);
and (n1266, n1262_mux, n1265_mux);
and (n1267, n385_mux, n322_mux);
not(n1268, n322_mux);
nor (n1269, n1267_mux, n1268_mux);
and (n1270, n1265_mux, n1269_mux);
and (n1271, n1262_mux, n1269_mux);
or (n1272_1, n1270_mux, n1271_mux);
or (n1272, n1266_mux, n1272_1);
and (n347, n325_mux, n319_mux);
and (n348, n334_mux, n322_mux);
and (n362, n347_mux, n348_mux);
buf(n42, g23_mux);
buf(n326, n42_mux);
and (n351, n350_mux, n326_mux);
and (n363, n348_mux, n351_mux);
and (n364, n347_mux, n351_mux);
or (n365_1, n363_mux, n364_mux);
or (n365, n362_mux, n365_1);
xor (n368, n366_mux, n367_mux);
xor (n370, n368_mux, n369_mux);
and (n1273, n365_mux, n370_mux);
xor (n374, n372_mux, n373_mux);
xor (n376, n374_mux, n375_mux);
and (n1274, n370_mux, n376_mux);
and (n1275, n365_mux, n376_mux);
or (n1276_1, n1274_mux, n1275_mux);
or (n1276, n1273_mux, n1276_1);
xor (n1277, n1262_mux, n1265_mux);
xor (n1278, n1277_mux, n1269_mux);
and (n1279, n1276_mux, n1278_mux);
xor (n1280, n1233_mux, n1235_mux);
xor (n1281, n1280_mux, n1237_mux);
and (n1282, n1278_mux, n1281_mux);
and (n1283, n1276_mux, n1281_mux);
or (n1284_1, n1282_mux, n1283_mux);
or (n1284, n1279_mux, n1284_1);
and (n1285, n1272_mux, n1284_mux);
xor (n1286, n1240_mux, n1242_mux);
xor (n1287, n1286_mux, n1245_mux);
and (n1288, n1284_mux, n1287_mux);
and (n1289, n1272_mux, n1287_mux);
or (n1290_1, n1288_mux, n1289_mux);
or (n1290, n1285_mux, n1290_1);
and (n1291, n1258_mux, n1290_mux);
xor (n1292, n1258_mux, n1290_mux);
xor (n1293, n1272_mux, n1284_mux);
xor (n1294, n1293_mux, n1287_mux);
buf(g356, g7_mux);
buf(n306, g356_mux);
not(n379, n306_mux);
and (n382, n381_mux, n306_mux);
nor (n383, n379_mux, n382_mux);
and (n386, n385_mux, n326_mux);
not(n387, n326_mux);
nor (n388, n386_mux, n387_mux);
and (n1295, n383_mux, n388_mux);
and (n333, n325_mux, n322_mux);
and (n335, n334_mux, n326_mux);
and (n343, n333_mux, n335_mux);
and (n345, n321_mux, n344_mux);
and (n358, n343_mux, n345_mux);
xor (n349, n347_mux, n348_mux);
xor (n352, n349_mux, n351_mux);
and (n359, n345_mux, n352_mux);
and (n360, n343_mux, n352_mux);
or (n361_1, n359_mux, n360_mux);
or (n361, n358_mux, n361_1);
xor (n371, n365_mux, n370_mux);
xor (n377, n371_mux, n376_mux);
and (n1296, n361_mux, n377_mux);
xor (n389, n383_mux, n388_mux);
and (n1297, n377_mux, n389_mux);
and (n1298, n361_mux, n389_mux);
or (n1299_1, n1297_mux, n1298_mux);
or (n1299, n1296_mux, n1299_1);
and (n1300, n1295_mux, n1299_mux);
xor (n1301, n1276_mux, n1278_mux);
xor (n1302, n1301_mux, n1281_mux);
and (n1303, n1299_mux, n1302_mux);
and (n1304, n1295_mux, n1302_mux);
or (n1305_1, n1303_mux, n1304_mux);
or (n1305, n1300_mux, n1305_1);
and (n1306, n1294_mux, n1305_mux);
xor (n1307, n1294_mux, n1305_mux);
xor (n1308, n1295_mux, n1299_mux);
xor (n1309, n1308_mux, n1302_mux);
and (n308, n306_mux, n307_mux);
and (n311, n309_mux, n310_mux);
and (n312, n308_mux, n311_mux);
and (n315, n313_mux, n314_mux);
and (n316, n311_mux, n315_mux);
and (n317, n308_mux, n315_mux);
or (n318_1, n316_mux, n317_mux);
or (n318, n312_mux, n318_1);
and (n320, n313_mux, n319_mux);
and (n323, n321_mux, n322_mux);
and (n324, n320_mux, n323_mux);
and (n327, n325_mux, n326_mux);
and (n328, n323_mux, n327_mux);
and (n329, n320_mux, n327_mux);
or (n330_1, n328_mux, n329_mux);
or (n330, n324_mux, n330_1);
and (n331, n321_mux, n319_mux);
and (n332, n330_mux, n331_mux);
xor (n336, n333_mux, n335_mux);
and (n337, n331_mux, n336_mux);
and (n338, n330_mux, n336_mux);
or (n339_1, n337_mux, n338_mux);
or (n339, n332_mux, n339_1);
xor (n340, n308_mux, n311_mux);
xor (n341, n340_mux, n315_mux);
and (n342, n339_mux, n341_mux);
xor (n346, n343_mux, n345_mux);
xor (n353, n346_mux, n352_mux);
and (n354, n341_mux, n353_mux);
and (n355, n339_mux, n353_mux);
or (n356_1, n354_mux, n355_mux);
or (n356, n342_mux, n356_1);
and (n1310, n318_mux, n356_mux);
xor (n378, n361_mux, n377_mux);
xor (n390, n378_mux, n389_mux);
and (n1311, n356_mux, n390_mux);
and (n1312, n318_mux, n390_mux);
or (n1313_1, n1311_mux, n1312_mux);
or (n1313, n1310_mux, n1313_1);
and (n1314, n1309_mux, n1313_mux);
xor (n1315, n1309_mux, n1313_mux);
xor (n357, n318_mux, n356_mux);
xor (n391, n357_mux, n390_mux);
and (n392, n309_mux, n314_mux);
and (n393, n313_mux, n344_mux);
and (n394, n392_mux, n393_mux);
and (n395, n309_mux, n319_mux);
and (n396, n313_mux, n322_mux);
and (n397, n395_mux, n396_mux);
and (n398, n321_mux, n326_mux);
and (n399, n396_mux, n398_mux);
and (n400, n395_mux, n398_mux);
or (n401_1, n399_mux, n400_mux);
or (n401, n397_mux, n401_1);
and (n402, n309_mux, n344_mux);
and (n403, n401_mux, n402_mux);
xor (n404, n320_mux, n323_mux);
xor (n405, n404_mux, n327_mux);
and (n406, n402_mux, n405_mux);
and (n407, n401_mux, n405_mux);
or (n408_1, n406_mux, n407_mux);
or (n408, n403_mux, n408_1);
xor (n409, n392_mux, n393_mux);
and (n410, n408_mux, n409_mux);
xor (n411, n330_mux, n331_mux);
xor (n412, n411_mux, n336_mux);
and (n413, n409_mux, n412_mux);
and (n414, n408_mux, n412_mux);
or (n415_1, n413_mux, n414_mux);
or (n415, n410_mux, n415_1);
and (n416, n394_mux, n415_mux);
xor (n417, n339_mux, n341_mux);
xor (n418, n417_mux, n353_mux);
and (n419, n415_mux, n418_mux);
and (n420, n394_mux, n418_mux);
or (n421_1, n419_mux, n420_mux);
or (n421, n416_mux, n421_1);
and (n1316, n391_mux, n421_mux);
xor (n422, n391_mux, n421_mux);
xor (n423, n394_mux, n415_mux);
xor (n424, n423_mux, n418_mux);
and (n425, n306_mux, n319_mux);
and (n426, n309_mux, n322_mux);
and (n427, n425_mux, n426_mux);
and (n428, n313_mux, n326_mux);
and (n429, n426_mux, n428_mux);
and (n430, n425_mux, n428_mux);
or (n431_1, n429_mux, n430_mux);
or (n431, n427_mux, n431_1);
and (n432, n306_mux, n344_mux);
and (n433, n431_mux, n432_mux);
xor (n434, n395_mux, n396_mux);
xor (n435, n434_mux, n398_mux);
and (n436, n432_mux, n435_mux);
and (n437, n431_mux, n435_mux);
or (n438_1, n436_mux, n437_mux);
or (n438, n433_mux, n438_1);
and (n439, n306_mux, n314_mux);
and (n440, n438_mux, n439_mux);
xor (n441, n401_mux, n402_mux);
xor (n442, n441_mux, n405_mux);
and (n443, n439_mux, n442_mux);
and (n444, n438_mux, n442_mux);
or (n445_1, n443_mux, n444_mux);
or (n445, n440_mux, n445_1);
xor (n446, n408_mux, n409_mux);
xor (n447, n446_mux, n412_mux);
and (n448, n445_mux, n447_mux);
and (n449, n424_mux, n448_mux);
xor (n450, n424_mux, n448_mux);
and (n451, n306_mux, n310_mux);
xor (n452, n445_mux, n447_mux);
and (n453, n451_mux, n452_mux);
xor (n454, n451_mux, n452_mux);
xor (n455, n438_mux, n439_mux);
xor (n456, n455_mux, n442_mux);
xor (n457, n431_mux, n432_mux);
xor (n458, n457_mux, n435_mux);
xor (n459, n425_mux, n426_mux);
xor (n460, n459_mux, n428_mux);
and (n461, n306_mux, n322_mux);
and (n462, n309_mux, n326_mux);
and (n463, n461_mux, n462_mux);
and (n464, n460_mux, n463_mux);
and (n465, n458_mux, n464_mux);
and (n466, n456_mux, n465_mux);
and (n467, n454_mux, n466_mux);
or (n468, n453_mux, n467_mux);
and (n469, n450_mux, n468_mux);
or (n470, n449_mux, n469_mux);
and (n1317, n422_mux, n470_mux);
or (n1318, n1316_mux, n1317_mux);
and (n1319, n1315_mux, n1318_mux);
or (n1320, n1314_mux, n1319_mux);
and (n1321, n1307_mux, n1320_mux);
or (n1322, n1306_mux, n1321_mux);
and (n1323, n1292_mux, n1322_mux);
or (n1324, n1291_mux, n1323_mux);
and (n1325, n1256_mux, n1324_mux);
or (n1326, n1255_mux, n1325_mux);
and (n1327, n1216_mux, n1326_mux);
or (n1328, n1215_mux, n1327_mux);
and (n1329, n1179_mux, n1328_mux);
or (n1330, n1178_mux, n1329_mux);
and (n1331, n1136_mux, n1330_mux);
or (n1332, n1135_mux, n1331_mux);
buf(n1333, n1332_mux);
buf(n1463, n1333_mux);
xor (n1334, n1136_mux, n1330_mux);
buf(n1335, n1334_mux);
buf(n1464, n1335_mux);
xor (n1336, n1179_mux, n1328_mux);
buf(n1337, n1336_mux);
buf(n1465, n1337_mux);
xor (n1338, n1216_mux, n1326_mux);
buf(n1339, n1338_mux);
buf(n1466, n1339_mux);
xor (n1340, n1256_mux, n1324_mux);
buf(n1341, n1340_mux);
buf(n1467, n1341_mux);
xor (n1342, n1292_mux, n1322_mux);
buf(n1343, n1342_mux);
buf(n1468, n1343_mux);
xor (n1344, n1307_mux, n1320_mux);
buf(n1345, n1344_mux);
buf(n1469, n1345_mux);
xor (n638, n450_mux, n468_mux);
buf(n639, n638_mux);
buf(n640, n639_mux);
buf(n33, g14_mux);
buf(n474, n33_mux);
buf(n46, g27_mux);
buf(n479, n46_mux);
and (n557, n474_mux, n479_mux);
buf(n32, g13_mux);
buf(n478, n32_mux);
buf(n47, g28_mux);
buf(n509, n47_mux);
and (n558, n478_mux, n509_mux);
and (n559, n557_mux, n558_mux);
buf(n48, g29_mux);
buf(n484, n48_mux);
and (n560, n474_mux, n484_mux);
buf(n49, g30_mux);
buf(n487, n49_mux);
and (n561, n478_mux, n487_mux);
and (n562, n560_mux, n561_mux);
buf(n31, g12_mux);
buf(n486, n31_mux);
buf(n50, g31_mux);
buf(n491, n50_mux);
and (n563, n486_mux, n491_mux);
and (n564, n561_mux, n563_mux);
and (n565, n560_mux, n563_mux);
or (n566_1, n564_mux, n565_mux);
or (n566, n562_mux, n566_1);
and (n567, n474_mux, n509_mux);
and (n568, n566_mux, n567_mux);
and (n485, n478_mux, n484_mux);
and (n488, n486_mux, n487_mux);
xor (n569, n485_mux, n488_mux);
buf(n30, g11_mux);
buf(n490, n30_mux);
and (n492, n490_mux, n491_mux);
xor (n570, n569_mux, n492_mux);
and (n571, n567_mux, n570_mux);
and (n572, n566_mux, n570_mux);
or (n573_1, n571_mux, n572_mux);
or (n573, n568_mux, n573_1);
xor (n574, n557_mux, n558_mux);
and (n575, n573_mux, n574_mux);
and (n489, n485_mux, n488_mux);
and (n493, n488_mux, n492_mux);
and (n494, n485_mux, n492_mux);
or (n495_1, n493_mux, n494_mux);
or (n495, n489_mux, n495_1);
and (n496, n486_mux, n484_mux);
xor (n576, n495_mux, n496_mux);
and (n498, n490_mux, n487_mux);
buf(n29, g10_mux);
buf(n499, n29_mux);
and (n500, n499_mux, n491_mux);
xor (n501, n498_mux, n500_mux);
xor (n577, n576_mux, n501_mux);
and (n578, n574_mux, n577_mux);
and (n579, n573_mux, n577_mux);
or (n580_1, n578_mux, n579_mux);
or (n580, n575_mux, n580_1);
xor (n588, n559_mux, n580_mux);
and (n497, n495_mux, n496_mux);
and (n502, n496_mux, n501_mux);
and (n503, n495_mux, n501_mux);
or (n504_1, n502_mux, n503_mux);
or (n504, n497_mux, n504_1);
buf(n34, g15_mux);
buf(n471, n34_mux);
buf(n44, g25_mux);
buf(n472, n44_mux);
and (n473, n471_mux, n472_mux);
buf(n45, g26_mux);
buf(n475, n45_mux);
and (n476, n474_mux, n475_mux);
xor (n505, n473_mux, n476_mux);
and (n480, n478_mux, n479_mux);
xor (n506, n505_mux, n480_mux);
xor (n582, n504_mux, n506_mux);
and (n508, n498_mux, n500_mux);
and (n510, n486_mux, n509_mux);
xor (n511, n508_mux, n510_mux);
and (n512, n490_mux, n484_mux);
and (n513, n499_mux, n487_mux);
xor (n514, n512_mux, n513_mux);
buf(n28, g9_mux);
buf(n515, n28_mux);
and (n516, n515_mux, n491_mux);
xor (n517, n514_mux, n516_mux);
xor (n518, n511_mux, n517_mux);
xor (n583, n582_mux, n518_mux);
xor (n589, n588_mux, n583_mux);
and (n590, n471_mux, n484_mux);
and (n591, n474_mux, n487_mux);
and (n592, n590_mux, n591_mux);
and (n593, n478_mux, n491_mux);
and (n594, n591_mux, n593_mux);
and (n595, n590_mux, n593_mux);
or (n596_1, n594_mux, n595_mux);
or (n596, n592_mux, n596_1);
and (n597, n471_mux, n509_mux);
and (n598, n596_mux, n597_mux);
xor (n599, n560_mux, n561_mux);
xor (n600, n599_mux, n563_mux);
and (n601, n597_mux, n600_mux);
and (n602, n596_mux, n600_mux);
or (n603_1, n601_mux, n602_mux);
or (n603, n598_mux, n603_1);
and (n604, n471_mux, n479_mux);
and (n605, n603_mux, n604_mux);
xor (n606, n566_mux, n567_mux);
xor (n607, n606_mux, n570_mux);
and (n608, n604_mux, n607_mux);
and (n609, n603_mux, n607_mux);
or (n610_1, n608_mux, n609_mux);
or (n610, n605_mux, n610_1);
xor (n611, n573_mux, n574_mux);
xor (n612, n611_mux, n577_mux);
and (n613, n610_mux, n612_mux);
xor (n615, n589_mux, n613_mux);
and (n616, n471_mux, n475_mux);
xor (n617, n610_mux, n612_mux);
and (n618, n616_mux, n617_mux);
xor (n619, n616_mux, n617_mux);
xor (n620, n603_mux, n604_mux);
xor (n621, n620_mux, n607_mux);
xor (n622, n596_mux, n597_mux);
xor (n623, n622_mux, n600_mux);
xor (n624, n590_mux, n591_mux);
xor (n625, n624_mux, n593_mux);
and (n626, n471_mux, n487_mux);
and (n627, n474_mux, n491_mux);
and (n628, n626_mux, n627_mux);
and (n629, n625_mux, n628_mux);
and (n630, n623_mux, n629_mux);
and (n631, n621_mux, n630_mux);
and (n632, n619_mux, n631_mux);
or (n633, n618_mux, n632_mux);
xor (n641, n615_mux, n633_mux);
buf(n642, n641_mux);
buf(n643, n642_mux);
and (n644, n640_mux, n643_mux);
xor (n645, n454_mux, n466_mux);
buf(n646, n645_mux);
buf(n647, n646_mux);
xor (n648, n619_mux, n631_mux);
buf(n649, n648_mux);
buf(n650, n649_mux);
and (n651, n647_mux, n650_mux);
xor (n652, n456_mux, n465_mux);
buf(n653, n652_mux);
buf(n654, n653_mux);
xor (n655, n621_mux, n630_mux);
buf(n656, n655_mux);
buf(n657, n656_mux);
and (n658, n654_mux, n657_mux);
xor (n659, n458_mux, n464_mux);
buf(n660, n659_mux);
buf(n661, n660_mux);
xor (n662, n623_mux, n629_mux);
buf(n663, n662_mux);
buf(n664, n663_mux);
and (n665, n661_mux, n664_mux);
xor (n666, n460_mux, n463_mux);
buf(n667, n666_mux);
buf(n668, n667_mux);
xor (n669, n625_mux, n628_mux);
buf(n670, n669_mux);
buf(n671, n670_mux);
and (n672, n668_mux, n671_mux);
xor (n673, n461_mux, n462_mux);
buf(n674, n673_mux);
buf(n675, n674_mux);
xor (n676, n626_mux, n627_mux);
buf(n677, n676_mux);
buf(n678, n677_mux);
and (n679, n675_mux, n678_mux);
and (n680, n306_mux, n326_mux);
buf(n681, n680_mux);
buf(n682, n681_mux);
and (n683, n471_mux, n491_mux);
buf(n684, n683_mux);
buf(n685, n684_mux);
and (n686, n682_mux, n685_mux);
and (n687, n678_mux, n686_mux);
and (n688, n675_mux, n686_mux);
or (n689_1, n687_mux, n688_mux);
or (n689, n679_mux, n689_1);
and (n690, n671_mux, n689_mux);
and (n691, n668_mux, n689_mux);
or (n692_1, n690_mux, n691_mux);
or (n692, n672_mux, n692_1);
and (n693, n664_mux, n692_mux);
and (n694, n661_mux, n692_mux);
or (n695_1, n693_mux, n694_mux);
or (n695, n665_mux, n695_1);
and (n696, n657_mux, n695_mux);
and (n697, n654_mux, n695_mux);
or (n698_1, n696_mux, n697_mux);
or (n698, n658_mux, n698_1);
and (n699, n650_mux, n698_mux);
and (n700, n647_mux, n698_mux);
or (n701_1, n699_mux, n700_mux);
or (n701, n651_mux, n701_1);
and (n702, n643_mux, n701_mux);
and (n703, n640_mux, n701_mux);
or (n704_1, n702_mux, n703_mux);
or (n704, n644_mux, n704_1);
xor (n705, t_0, n704_mux);
buf(n706, n705_mux);
not(n25, n706_mux);
buf(n816, n35_mux);
buf(n43, g24_mux);
buf(n817, n43_mux);
and (n835, n816_mux, n817_mux);
buf(n797, n36_mux);
buf(n798, n44_mux);
and (n819, n797_mux, n798_mux);
buf(n778, n37_mux);
buf(n779, n45_mux);
and (n800, n778_mux, n779_mux);
buf(n759, n38_mux);
buf(n760, n46_mux);
and (n781, n759_mux, n760_mux);
buf(n740, n39_mux);
buf(n741, n47_mux);
and (n762, n740_mux, n741_mux);
buf(n721, n40_mux);
buf(n722, n48_mux);
and (n743, n721_mux, n722_mux);
buf(n708, n41_mux);
buf(n709, n49_mux);
and (n724, n708_mux, n709_mux);
buf(n298, n42_mux);
buf(n299, n50_mux);
and (n711, n298_mux, n299_mux);
and (n725, n709_mux, n711_mux);
and (n726, n708_mux, n711_mux);
or (n727_1, n725_mux, n726_mux);
or (n727, n724_mux, n727_1);
and (n744, n722_mux, n727_mux);
and (n745, n721_mux, n727_mux);
or (n746_1, n744_mux, n745_mux);
or (n746, n743_mux, n746_1);
and (n763, n741_mux, n746_mux);
and (n764, n740_mux, n746_mux);
or (n765_1, n763_mux, n764_mux);
or (n765, n762_mux, n765_1);
and (n782, n760_mux, n765_mux);
and (n783, n759_mux, n765_mux);
or (n784_1, n782_mux, n783_mux);
or (n784, n781_mux, n784_1);
and (n801, n779_mux, n784_mux);
and (n802, n778_mux, n784_mux);
or (n803_1, n801_mux, n802_mux);
or (n803, n800_mux, n803_1);
and (n820, n798_mux, n803_mux);
and (n821, n797_mux, n803_mux);
or (n822_1, n820_mux, n821_mux);
or (n822, n819_mux, n822_1);
and (n836, n817_mux, n822_mux);
and (n837, n816_mux, n822_mux);
or (n838_1, n836_mux, n837_mux);
or (n838, n835_mux, n838_1);
buf(n839, n838_mux);
and (n26, n25_mux, n839_mux);
buf(n825, g349_mux);
buf(g357, g8_mux);
buf(n826, g357_mux);
and (n840, n825_mux, n826_mux);
buf(n806, g350_mux);
buf(n807, n28_mux);
and (n828, n806_mux, n807_mux);
buf(n787, g351_mux);
buf(n788, n29_mux);
and (n809, n787_mux, n788_mux);
buf(n768, g352_mux);
buf(n769, n30_mux);
and (n790, n768_mux, n769_mux);
buf(n749, g353_mux);
buf(n750, n31_mux);
and (n771, n749_mux, n750_mux);
buf(n730, g354_mux);
buf(n731, n32_mux);
and (n752, n730_mux, n731_mux);
buf(n714, g355_mux);
buf(n715, n33_mux);
and (n733, n714_mux, n715_mux);
buf(n302, g356_mux);
buf(n303, n34_mux);
and (n717, n302_mux, n303_mux);
and (n734, n715_mux, n717_mux);
and (n735, n714_mux, n717_mux);
or (n736_1, n734_mux, n735_mux);
or (n736, n733_mux, n736_1);
and (n753, n731_mux, n736_mux);
and (n754, n730_mux, n736_mux);
or (n755_1, n753_mux, n754_mux);
or (n755, n752_mux, n755_1);
and (n772, n750_mux, n755_mux);
and (n773, n749_mux, n755_mux);
or (n774_1, n772_mux, n773_mux);
or (n774, n771_mux, n774_1);
and (n791, n769_mux, n774_mux);
and (n792, n768_mux, n774_mux);
or (n793_1, n791_mux, n792_mux);
or (n793, n790_mux, n793_1);
and (n810, n788_mux, n793_mux);
and (n811, n787_mux, n793_mux);
or (n812_1, n810_mux, n811_mux);
or (n812, n809_mux, n812_1);
and (n829, n807_mux, n812_mux);
and (n830, n806_mux, n812_mux);
or (n831_1, n829_mux, n830_mux);
or (n831, n828_mux, n831_1);
and (n841, n826_mux, n831_mux);
and (n842, n825_mux, n831_mux);
or (n843_1, n841_mux, n842_mux);
or (n843, n840_mux, n843_1);
buf(n844, n843_mux);
and (n27, n844_mux, n706_mux);
or (n845, n26_mux, n27_mux);
buf(n1454, n845_mux);
xor (n1346, n1315_mux, n1318_mux);
buf(n1347, n1346_mux);
buf(n1470, n1347_mux);
and (n1478, n1454_mux, n1470_mux);
not(n22, n706_mux);
xor (n818, n816_mux, n817_mux);
xor (n823, n818_mux, n822_mux);
buf(n824, n823_mux);
and (n23, n22_mux, n824_mux);
xor (n827, n825_mux, n826_mux);
xor (n832, n827_mux, n831_mux);
buf(n833, n832_mux);
and (n24, n833_mux, n706_mux);
or (n834, n23_mux, n24_mux);
buf(n1455, n834_mux);
and (n1479, n1455_mux, t_1);
not(n19, n706_mux);
xor (n799, n797_mux, n798_mux);
xor (n804, n799_mux, n803_mux);
buf(n805, n804_mux);
and (n20, n19_mux, n805_mux);
xor (n808, n806_mux, n807_mux);
xor (n813, n808_mux, n812_mux);
buf(n814, n813_mux);
and (n21, n814_mux, n706_mux);
or (n815, n20_mux, n21_mux);
buf(n1456, n815_mux);
buf(n1471, n639_mux);
and (n1480, n1456_mux, n1471_mux);
not(n16, n706_mux);
xor (n780, n778_mux, n779_mux);
xor (n785, n780_mux, n784_mux);
buf(n786, n785_mux);
and (n17, n16_mux, n786_mux);
xor (n789, n787_mux, n788_mux);
xor (n794, n789_mux, n793_mux);
buf(n795, n794_mux);
and (n18, n795_mux, n706_mux);
or (n796, n17_mux, n18_mux);
buf(n1457, n796_mux);
buf(n1472, n646_mux);
and (n1481, n1457_mux, n1472_mux);
not(n13, n706_mux);
xor (n761, n759_mux, n760_mux);
xor (n766, n761_mux, n765_mux);
buf(n767, n766_mux);
and (n14, n13_mux, n767_mux);
xor (n770, n768_mux, n769_mux);
xor (n775, n770_mux, n774_mux);
buf(n776, n775_mux);
and (n15, n776_mux, n706_mux);
or (n777, n14_mux, n15_mux);
buf(n1458, n777_mux);
buf(n1473, n653_mux);
and (n1482, n1458_mux, n1473_mux);
not(n10, n706_mux);
xor (n742, n740_mux, n741_mux);
xor (n747, n742_mux, n746_mux);
buf(n748, n747_mux);
and (n11, n10_mux, n748_mux);
xor (n751, n749_mux, n750_mux);
xor (n756, n751_mux, n755_mux);
buf(n757, n756_mux);
and (n12, n757_mux, n706_mux);
or (n758, n11_mux, n12_mux);
buf(n1459, n758_mux);
buf(n1474, n660_mux);
and (n1483, n1459_mux, n1474_mux);
not(n7, n706_mux);
xor (n723, n721_mux, n722_mux);
xor (n728, n723_mux, n727_mux);
buf(n729, n728_mux);
and (n8, n7_mux, n729_mux);
xor (n732, n730_mux, n731_mux);
xor (n737, n732_mux, n736_mux);
buf(n738, n737_mux);
and (n9, n738_mux, n706_mux);
or (n739, n8_mux, n9_mux);
buf(n1460, n739_mux);
buf(n1475, n667_mux);
and (n1484, n1460_mux, n1475_mux);
not(n4, n706_mux);
xor (n710, n708_mux, n709_mux);
xor (n712, n710_mux, n711_mux);
buf(n713, n712_mux);
and (n5, n4_mux, n713_mux);
xor (n716, n714_mux, n715_mux);
xor (n718, n716_mux, n717_mux);
buf(n719, n718_mux);
and (n6, n719_mux, n706_mux);
or (n720, n5_mux, n6_mux);
buf(n1461, n720_mux);
buf(n1476, n674_mux);
and (n1485, n1461_mux, n1476_mux);
not(n1, n706_mux);
xor (n300, n298_mux, n299_mux);
buf(n301, n300_mux);
and (n2, n1_mux, n301_mux);
xor (n304, n302_mux, n303_mux);
buf(n305, n304_mux);
and (n3, n305_mux, n706_mux);
or (n707, n2_mux, n3_mux);
buf(n1462, n707_mux);
buf(n1477, n681_mux);
and (n1486, n1462_mux, n1477_mux);
and (n1487, n1476_mux, n1486_mux);
and (n1488, n1461_mux, n1486_mux);
or (n1489_1, n1487_mux, n1488_mux);
or (n1489, n1485_mux, n1489_1);
and (n1490, n1475_mux, n1489_mux);
and (n1491, n1460_mux, n1489_mux);
or (n1492_1, n1490_mux, n1491_mux);
or (n1492, n1484_mux, n1492_1);
and (n1493, n1474_mux, n1492_mux);
and (n1494, n1459_mux, n1492_mux);
or (n1495_1, n1493_mux, n1494_mux);
or (n1495, n1483_mux, n1495_1);
and (n1496, n1473_mux, n1495_mux);
and (n1497, n1458_mux, n1495_mux);
or (n1498_1, n1496_mux, n1497_mux);
or (n1498, n1482_mux, n1498_1);
and (n1499, n1472_mux, n1498_mux);
and (n1500, n1457_mux, n1498_mux);
or (n1501_1, n1499_mux, n1500_mux);
or (n1501, n1481_mux, n1501_1);
and (n1502, n1471_mux, n1501_mux);
and (n1503, n1456_mux, n1501_mux);
or (n1504_1, n1502_mux, n1503_mux);
or (n1504, n1480_mux, n1504_1);
and (n1505, t_1, n1504_mux);
and (n1506, n1455_mux, n1504_mux);
or (n1507_1, n1505_mux, n1506_mux);
or (n1507, n1479_mux, n1507_1);
and (n1508, n1470_mux, n1507_mux);
and (n1509, n1454_mux, n1507_mux);
or (n1510_1, n1508_mux, n1509_mux);
or (n1510, n1478_mux, n1510_1);
and (n1511, n1469_mux, n1510_mux);
and (n1512, n1468_mux, n1511_mux);
and (n1513, n1467_mux, n1512_mux);
and (n1514, n1466_mux, n1513_mux);
and (n1515, n1465_mux, n1514_mux);
and (n1516, n1464_mux, n1515_mux);
and (n1517, n1463_mux, n1516_mux);
buf(n1518, n1517_mux);
buf(n99, n1518_mux);
buf(g80, n99);
xor (n1519, n1463_mux, n1516_mux);
buf(n1520, n1519_mux);
buf(n100, n1520_mux);
buf(g81, n100);
xor (n1521, n1464_mux, n1515_mux);
buf(n1522, n1521_mux);
buf(n101, n1522_mux);
buf(g82, n101);
xor (n1523, n1465_mux, n1514_mux);
buf(n1524, n1523_mux);
buf(n102, n1524_mux);
buf(g83, n102);
xor (n1525, n1466_mux, n1513_mux);
buf(n1526, n1525_mux);
buf(n103, n1526_mux);
buf(g84, n103);
xor (n1527, n1467_mux, n1512_mux);
buf(n1528, n1527_mux);
buf(n104, n1528_mux);
buf(g85, n104);
xor (n1529, n1468_mux, n1511_mux);
buf(n1530, n1529_mux);
buf(n105, n1530_mux);
buf(g86, n105);
xor (n1531, n1469_mux, n1510_mux);
buf(n1532, n1531_mux);
buf(n106, n1532_mux);
buf(g87, n106);
xor (n1533, n1454_mux, n1470_mux);
xor (n1534, n1533_mux, n1507_mux);
buf(n1535, n1534_mux);
buf(n107, n1535_mux);
buf(g88, n107);
xor (n1536, n1455_mux, t_1);
xor (n1537, n1536_mux, n1504_mux);
buf(n1538, n1537_mux);
buf(n108, n1538_mux);
buf(g89, n108);
xor (n1539, n1456_mux, n1471_mux);
xor (n1540, n1539_mux, n1501_mux);
buf(n1541, n1540_mux);
buf(n109, n1541_mux);
buf(g90, n109);
xor (n1542, n1457_mux, n1472_mux);
xor (n1543, n1542_mux, n1498_mux);
buf(n1544, n1543_mux);
buf(n110, n1544_mux);
buf(g91, n110);
xor (n1545, n1458_mux, n1473_mux);
xor (n1546, n1545_mux, n1495_mux);
buf(n1547, n1546_mux);
buf(n111, n1547_mux);
buf(g92, n111);
xor (n1548, n1459_mux, n1474_mux);
xor (n1549, n1548_mux, n1492_mux);
buf(n1550, n1549_mux);
buf(n112, n1550_mux);
buf(g93, n112);
xor (n1551, n1460_mux, n1475_mux);
xor (n1552, n1551_mux, n1489_mux);
buf(n1553, n1552_mux);
buf(n113, n1553_mux);
buf(g94, n113);
xor (n1554, n1461_mux, n1476_mux);
xor (n1555, n1554_mux, n1486_mux);
buf(n1556, n1555_mux);
buf(n114, n1556_mux);
buf(g95, n114);
xor (n1557, n1462_mux, n1477_mux);
buf(n1558, n1557_mux);
buf(n115, n1558_mux);
buf(g96, n115);
buf(n116, 1'b0);
buf(g97, n116);
buf(n117, 1'b0);
buf(g98, n117);
buf(n118, 1'b0);
buf(g99, n118);
buf(n119, 1'b0);
buf(g100, n119);
buf(n120, 1'b0);
buf(g101, n120);
buf(n121, 1'b0);
buf(g102, n121);
buf(n122, 1'b0);
buf(g103, n122);
buf(n123, 1'b0);
buf(g104, n123);
buf(n124, 1'b0);
buf(g105, n124);
buf(n125, 1'b0);
buf(g106, n125);
buf(n126, 1'b0);
buf(g107, n126);
buf(n127, 1'b0);
buf(g108, n127);
buf(n128, 1'b0);
buf(g109, n128);
buf(n129, 1'b0);
buf(g110, n129);
buf(n130, 1'b0);
buf(g111, n130);
buf(n131, 1'b0);
buf(g112, n131);
buf(n132, 1'b0);
buf(g113, n132);
buf(n133, 1'b0);
buf(g114, n133);
buf(n134, 1'b0);
buf(g115, n134);
buf(n135, 1'b0);
buf(g116, n135);
buf(n136, 1'b0);
buf(g117, n136);
buf(n137, 1'b0);
buf(g118, n137);
buf(n138, 1'b0);
buf(g119, n138);
buf(n139, 1'b0);
buf(g120, n139);
buf(n140, 1'b0);
buf(g121, n140);
buf(n141, 1'b0);
buf(g122, n141);
buf(n142, 1'b0);
buf(g123, n142);
buf(n143, 1'b0);
buf(g124, n143);
buf(n144, 1'b0);
buf(g125, n144);
buf(n145, 1'b0);
buf(g126, n145);
buf(n146, 1'b0);
buf(g127, n146);
buf(n147, 1'b0);
buf(g128, n147);
buf(n148, 1'b0);
buf(g129, n148);
buf(n149, 1'b0);
buf(g130, n149);
buf(n150, 1'b0);
buf(g131, n150);
buf(n151, 1'b0);
buf(g132, n151);
buf(n152, 1'b0);
buf(g133, n152);
buf(n153, 1'b0);
buf(g134, n153);
buf(n154, 1'b0);
buf(g135, n154);
buf(n155, 1'b0);
buf(g136, n155);
buf(n156, 1'b0);
buf(g137, n156);
buf(n157, 1'b0);
buf(g138, n157);
buf(n158, 1'b0);
buf(g139, n158);
buf(n159, 1'b0);
buf(g140, n159);
buf(n160, 1'b0);
buf(g141, n160);
buf(n161, 1'b0);
buf(g142, n161);
buf(n162, 1'b0);
buf(g143, n162);
buf(n549, g357_mux);
buf(n545, n43_mux);
and (n866, n549_mux, n545_mux);
not(n867, n490_mux);
not(n546, n545_mux);
and (n868, n546_mux, n490_mux);
nor (n869, n867_mux, n868_mux);
and (n870, n499_mux, n472_mux);
and (n871, n869_mux, n870_mux);
and (n872, n515_mux, n475_mux);
and (n873, n870_mux, n872_mux);
and (n874, n869_mux, n872_mux);
or (n875_1, n873_mux, n874_mux);
or (n875, n871_mux, n875_1);
not(n876, n499_mux);
and (n877, n546_mux, n499_mux);
nor (n878, n876_mux, n877_mux);
and (n879, n875_mux, n878_mux);
and (n880, n515_mux, n472_mux);
and (n881, n878_mux, n880_mux);
and (n882, n875_mux, n880_mux);
or (n883_1, n881_mux, n882_mux);
or (n883, n879_mux, n883_1);
not(n884, n515_mux);
and (n885, n546_mux, n515_mux);
nor (n886, n884_mux, n885_mux);
and (n887, n883_mux, n886_mux);
not(n550, n549_mux);
and (n888, n550_mux, n472_mux);
not(n889, n472_mux);
nor (n890, n888_mux, n889_mux);
and (n891, n886_mux, n890_mux);
and (n892, n883_mux, n890_mux);
or (n893_1, n891_mux, n892_mux);
or (n893, n887_mux, n893_1);
and (n894, n866_mux, n893_mux);
xor (n895, n866_mux, n893_mux);
xor (n896, n883_mux, n886_mux);
xor (n897, n896_mux, n890_mux);
not(n898, n486_mux);
and (n899, n546_mux, n486_mux);
nor (n900, n898_mux, n899_mux);
and (n901, n490_mux, n472_mux);
and (n902, n900_mux, n901_mux);
and (n903, n550_mux, n509_mux);
not(n904, n509_mux);
nor (n905, n903_mux, n904_mux);
and (n906, n901_mux, n905_mux);
and (n907, n900_mux, n905_mux);
or (n908_1, n906_mux, n907_mux);
or (n908, n902_mux, n908_1);
and (n909, n490_mux, n475_mux);
and (n910, n499_mux, n479_mux);
and (n911, n909_mux, n910_mux);
and (n912, n515_mux, n509_mux);
and (n913, n910_mux, n912_mux);
and (n914, n909_mux, n912_mux);
or (n915_1, n913_mux, n914_mux);
or (n915, n911_mux, n915_1);
and (n916, n499_mux, n475_mux);
and (n917, n915_mux, n916_mux);
and (n918, n515_mux, n479_mux);
and (n919, n916_mux, n918_mux);
and (n920, n915_mux, n918_mux);
or (n921_1, n919_mux, n920_mux);
or (n921, n917_mux, n921_1);
and (n922, n908_mux, n921_mux);
xor (n923, n869_mux, n870_mux);
xor (n924, n923_mux, n872_mux);
and (n925, n921_mux, n924_mux);
and (n926, n908_mux, n924_mux);
or (n927_1, n925_mux, n926_mux);
or (n927, n922_mux, n927_1);
and (n928, n550_mux, n475_mux);
not(n929, n475_mux);
nor (n930, n928_mux, n929_mux);
and (n931, n927_mux, n930_mux);
xor (n932, n875_mux, n878_mux);
xor (n933, n932_mux, n880_mux);
and (n934, n930_mux, n933_mux);
and (n935, n927_mux, n933_mux);
or (n936_1, n934_mux, n935_mux);
or (n936, n931_mux, n936_1);
and (n937, n897_mux, n936_mux);
xor (n938, n897_mux, n936_mux);
xor (n939, n927_mux, n930_mux);
xor (n940, n939_mux, n933_mux);
and (n941, n490_mux, n479_mux);
and (n942, n499_mux, n509_mux);
and (n943, n941_mux, n942_mux);
and (n944, n515_mux, n484_mux);
and (n945, n942_mux, n944_mux);
and (n946, n941_mux, n944_mux);
or (n947_1, n945_mux, n946_mux);
or (n947, n943_mux, n947_1);
and (n948, n478_mux, n472_mux);
and (n949, n486_mux, n475_mux);
and (n950, n948_mux, n949_mux);
and (n951, n947_mux, n950_mux);
xor (n952, n909_mux, n910_mux);
xor (n953, n952_mux, n912_mux);
and (n954, n950_mux, n953_mux);
and (n955, n947_mux, n953_mux);
or (n956_1, n954_mux, n955_mux);
or (n956, n951_mux, n956_1);
xor (n957, n900_mux, n901_mux);
xor (n958, n957_mux, n905_mux);
and (n959, n956_mux, n958_mux);
xor (n960, n915_mux, n916_mux);
xor (n961, n960_mux, n918_mux);
and (n962, n958_mux, n961_mux);
and (n963, n956_mux, n961_mux);
or (n964_1, n962_mux, n963_mux);
or (n964, n959_mux, n964_1);
and (n965, n550_mux, n479_mux);
not(n966, n479_mux);
nor (n967, n965_mux, n966_mux);
and (n968, n964_mux, n967_mux);
xor (n969, n908_mux, n921_mux);
xor (n970, n969_mux, n924_mux);
and (n971, n967_mux, n970_mux);
and (n972, n964_mux, n970_mux);
or (n973_1, n971_mux, n972_mux);
or (n973, n968_mux, n973_1);
and (n974, n940_mux, n973_mux);
xor (n975, n940_mux, n973_mux);
xor (n976, n964_mux, n967_mux);
xor (n977, n976_mux, n970_mux);
not(n978, n478_mux);
and (n979, n546_mux, n478_mux);
nor (n980, n978_mux, n979_mux);
and (n981, n486_mux, n472_mux);
and (n982, n980_mux, n981_mux);
and (n983, n550_mux, n484_mux);
not(n984, n484_mux);
nor (n985, n983_mux, n984_mux);
and (n986, n981_mux, n985_mux);
and (n987, n980_mux, n985_mux);
or (n988_1, n986_mux, n987_mux);
or (n988, n982_mux, n988_1);
and (n537, n490_mux, n509_mux);
and (n538, n499_mux, n484_mux);
and (n989, n537_mux, n538_mux);
and (n540, n515_mux, n487_mux);
and (n990, n538_mux, n540_mux);
and (n991, n537_mux, n540_mux);
or (n992_1, n990_mux, n991_mux);
or (n992, n989_mux, n992_1);
xor (n993, n941_mux, n942_mux);
xor (n994, n993_mux, n944_mux);
and (n995, n992_mux, n994_mux);
xor (n996, n948_mux, n949_mux);
and (n997, n994_mux, n996_mux);
and (n998, n992_mux, n996_mux);
or (n999_1, n997_mux, n998_mux);
or (n999, n995_mux, n999_1);
xor (n1000, n980_mux, n981_mux);
xor (n1001, n1000_mux, n985_mux);
and (n1002, n999_mux, n1001_mux);
xor (n1003, n947_mux, n950_mux);
xor (n1004, n1003_mux, n953_mux);
and (n1005, n1001_mux, n1004_mux);
and (n1006, n999_mux, n1004_mux);
or (n1007_1, n1005_mux, n1006_mux);
or (n1007, n1002_mux, n1007_1);
and (n1008, n988_mux, n1007_mux);
xor (n1009, n956_mux, n958_mux);
xor (n1010, n1009_mux, n961_mux);
and (n1011, n1007_mux, n1010_mux);
and (n1012, n988_mux, n1010_mux);
or (n1013_1, n1011_mux, n1012_mux);
or (n1013, n1008_mux, n1013_1);
and (n1014, n977_mux, n1013_mux);
xor (n1015, n977_mux, n1013_mux);
xor (n1016, n988_mux, n1007_mux);
xor (n1017, n1016_mux, n1010_mux);
and (n531, n474_mux, n472_mux);
and (n532, n478_mux, n475_mux);
and (n1018, n531_mux, n532_mux);
and (n534, n486_mux, n479_mux);
and (n1019, n532_mux, n534_mux);
and (n1020, n531_mux, n534_mux);
or (n1021_1, n1019_mux, n1020_mux);
or (n1021, n1018_mux, n1021_1);
not(n1022, n474_mux);
and (n1023, n546_mux, n474_mux);
nor (n1024, n1022_mux, n1023_mux);
and (n1025, n1021_mux, n1024_mux);
and (n1026, n550_mux, n487_mux);
not(n1027, n487_mux);
nor (n1028, n1026_mux, n1027_mux);
and (n1029, n1024_mux, n1028_mux);
and (n1030, n1021_mux, n1028_mux);
or (n1031_1, n1029_mux, n1030_mux);
or (n1031, n1025_mux, n1031_1);
and (n527, n512_mux, n513_mux);
and (n528, n513_mux, n516_mux);
and (n529, n512_mux, n516_mux);
or (n530_1, n528_mux, n529_mux);
or (n530, n527_mux, n530_1);
xor (n533, n531_mux, n532_mux);
xor (n535, n533_mux, n534_mux);
and (n1032, n530_mux, n535_mux);
xor (n539, n537_mux, n538_mux);
xor (n541, n539_mux, n540_mux);
and (n1033, n535_mux, n541_mux);
and (n1034, n530_mux, n541_mux);
or (n1035_1, n1033_mux, n1034_mux);
or (n1035, n1032_mux, n1035_1);
xor (n1036, n1021_mux, n1024_mux);
xor (n1037, n1036_mux, n1028_mux);
and (n1038, n1035_mux, n1037_mux);
xor (n1039, n992_mux, n994_mux);
xor (n1040, n1039_mux, n996_mux);
and (n1041, n1037_mux, n1040_mux);
and (n1042, n1035_mux, n1040_mux);
or (n1043_1, n1041_mux, n1042_mux);
or (n1043, n1038_mux, n1043_1);
and (n1044, n1031_mux, n1043_mux);
xor (n1045, n999_mux, n1001_mux);
xor (n1046, n1045_mux, n1004_mux);
and (n1047, n1043_mux, n1046_mux);
and (n1048, n1031_mux, n1046_mux);
or (n1049_1, n1047_mux, n1048_mux);
or (n1049, n1044_mux, n1049_1);
and (n1050, n1017_mux, n1049_mux);
xor (n1051, n1017_mux, n1049_mux);
xor (n1052, n1031_mux, n1043_mux);
xor (n1053, n1052_mux, n1046_mux);
not(n544, n471_mux);
and (n547, n546_mux, n471_mux);
nor (n548, n544_mux, n547_mux);
and (n551, n550_mux, n491_mux);
not(n552, n491_mux);
nor (n553, n551_mux, n552_mux);
and (n1054, n548_mux, n553_mux);
and (n523, n508_mux, n510_mux);
and (n524, n510_mux, n517_mux);
and (n525, n508_mux, n517_mux);
or (n526_1, n524_mux, n525_mux);
or (n526, n523_mux, n526_1);
xor (n536, n530_mux, n535_mux);
xor (n542, n536_mux, n541_mux);
and (n1055, n526_mux, n542_mux);
xor (n554, n548_mux, n553_mux);
and (n1056, n542_mux, n554_mux);
and (n1057, n526_mux, n554_mux);
or (n1058_1, n1056_mux, n1057_mux);
or (n1058, n1055_mux, n1058_1);
and (n1059, n1054_mux, n1058_mux);
xor (n1060, n1035_mux, n1037_mux);
xor (n1061, n1060_mux, n1040_mux);
and (n1062, n1058_mux, n1061_mux);
and (n1063, n1054_mux, n1061_mux);
or (n1064_1, n1062_mux, n1063_mux);
or (n1064, n1059_mux, n1064_1);
and (n1065, n1053_mux, n1064_mux);
xor (n1066, n1053_mux, n1064_mux);
xor (n1067, n1054_mux, n1058_mux);
xor (n1068, n1067_mux, n1061_mux);
and (n477, n473_mux, n476_mux);
and (n481, n476_mux, n480_mux);
and (n482, n473_mux, n480_mux);
or (n483_1, n481_mux, n482_mux);
or (n483, n477_mux, n483_1);
and (n507, n504_mux, n506_mux);
and (n519, n506_mux, n518_mux);
and (n520, n504_mux, n518_mux);
or (n521_1, n519_mux, n520_mux);
or (n521, n507_mux, n521_1);
and (n1069, n483_mux, n521_mux);
xor (n543, n526_mux, n542_mux);
xor (n555, n543_mux, n554_mux);
and (n1070, n521_mux, n555_mux);
and (n1071, n483_mux, n555_mux);
or (n1072_1, n1070_mux, n1071_mux);
or (n1072, n1069_mux, n1072_1);
and (n1073, n1068_mux, n1072_mux);
xor (n1074, n1068_mux, n1072_mux);
xor (n522, n483_mux, n521_mux);
xor (n556, n522_mux, n555_mux);
and (n581, n559_mux, n580_mux);
and (n584, n580_mux, n583_mux);
and (n585, n559_mux, n583_mux);
or (n586_1, n584_mux, n585_mux);
or (n586, n581_mux, n586_1);
and (n1075, n556_mux, n586_mux);
xor (n587, n556_mux, n586_mux);
and (n614, n589_mux, n613_mux);
and (n634, n615_mux, n633_mux);
or (n635, n614_mux, n634_mux);
and (n1076, n587_mux, n635_mux);
or (n1077, n1075_mux, n1076_mux);
and (n1078, n1074_mux, n1077_mux);
or (n1079, n1073_mux, n1078_mux);
and (n1080, n1066_mux, n1079_mux);
or (n1081, n1065_mux, n1080_mux);
and (n1082, n1051_mux, n1081_mux);
or (n1083, n1050_mux, n1082_mux);
and (n1084, n1015_mux, n1083_mux);
or (n1085, n1014_mux, n1084_mux);
and (n1086, n975_mux, n1085_mux);
or (n1087, n974_mux, n1086_mux);
and (n1088, n938_mux, n1087_mux);
or (n1089, n937_mux, n1088_mux);
and (n1090, n895_mux, n1089_mux);
or (n1091, n894_mux, n1090_mux);
buf(n1092, n1091_mux);
buf(n1357, n1092_mux);
xor (n1093, n895_mux, n1089_mux);
buf(n1094, n1093_mux);
buf(n1358, n1094_mux);
xor (n1095, n938_mux, n1087_mux);
buf(n1096, n1095_mux);
buf(n1359, n1096_mux);
xor (n1097, n975_mux, n1085_mux);
buf(n1098, n1097_mux);
buf(n1360, n1098_mux);
xor (n1099, n1015_mux, n1083_mux);
buf(n1100, n1099_mux);
buf(n1361, n1100_mux);
xor (n1101, n1051_mux, n1081_mux);
buf(n1102, n1101_mux);
buf(n1362, n1102_mux);
xor (n1103, n1066_mux, n1079_mux);
buf(n1104, n1103_mux);
buf(n1363, n1104_mux);
buf(n1348, n845_mux);
xor (n1105, n1074_mux, n1077_mux);
buf(n1106, n1105_mux);
buf(n1364, n1106_mux);
and (n1373, n1348_mux, n1364_mux);
buf(n1349, n834_mux);
xor (n636, n587_mux, n635_mux);
buf(n637, n636_mux);
buf(n1365, n637_mux);
and (n1374, n1349_mux, n1365_mux);
buf(n1350, n815_mux);
buf(n1366, n642_mux);
and (n1375, n1350_mux, n1366_mux);
buf(n1351, n796_mux);
buf(n1367, n649_mux);
and (n1376, n1351_mux, n1367_mux);
buf(n1352, n777_mux);
buf(n1368, n656_mux);
and (n1377, n1352_mux, n1368_mux);
buf(n1353, n758_mux);
buf(n1369, n663_mux);
and (n1378, n1353_mux, n1369_mux);
buf(n1354, n739_mux);
buf(n1370, n670_mux);
and (n1379, n1354_mux, n1370_mux);
buf(n1355, n720_mux);
buf(n1371, n677_mux);
and (n1380, n1355_mux, n1371_mux);
buf(n1356, n707_mux);
buf(n1372, n684_mux);
and (n1381, n1356_mux, n1372_mux);
and (n1382, n1371_mux, n1381_mux);
and (n1383, n1355_mux, n1381_mux);
or (n1384_1, n1382_mux, n1383_mux);
or (n1384, n1380_mux, n1384_1);
and (n1385, n1370_mux, n1384_mux);
and (n1386, n1354_mux, n1384_mux);
or (n1387_1, n1385_mux, n1386_mux);
or (n1387, n1379_mux, n1387_1);
and (n1388, n1369_mux, n1387_mux);
and (n1389, n1353_mux, n1387_mux);
or (n1390_1, n1388_mux, n1389_mux);
or (n1390, n1378_mux, n1390_1);
and (n1391, n1368_mux, n1390_mux);
and (n1392, n1352_mux, n1390_mux);
or (n1393_1, n1391_mux, n1392_mux);
or (n1393, n1377_mux, n1393_1);
and (n1394, n1367_mux, n1393_mux);
and (n1395, n1351_mux, n1393_mux);
or (n1396_1, n1394_mux, n1395_mux);
or (n1396, n1376_mux, n1396_1);
and (n1397, n1366_mux, n1396_mux);
and (n1398, n1350_mux, n1396_mux);
or (n1399_1, n1397_mux, n1398_mux);
or (n1399, n1375_mux, n1399_1);
and (n1400, n1365_mux, n1399_mux);
and (n1401, n1349_mux, n1399_mux);
or (n1402_1, n1400_mux, n1401_mux);
or (n1402, n1374_mux, n1402_1);
and (n1403, n1364_mux, n1402_mux);
and (n1404, n1348_mux, n1402_mux);
or (n1405_1, n1403_mux, n1404_mux);
or (n1405, n1373_mux, n1405_1);
and (n1406, n1363_mux, n1405_mux);
and (n1407, n1362_mux, n1406_mux);
and (n1408, n1361_mux, n1407_mux);
and (n1409, n1360_mux, n1408_mux);
and (n1410, n1359_mux, n1409_mux);
and (n1411, n1358_mux, n1410_mux);
and (n1412, n1357_mux, n1411_mux);
buf(n1413, n1412_mux);
buf(n163, n1413_mux);
buf(g144, n163);
xor (n1414, n1357_mux, n1411_mux);
buf(n1415, n1414_mux);
buf(n164, n1415_mux);
buf(g145, n164);
xor (n1416, n1358_mux, n1410_mux);
buf(n1417, n1416_mux);
buf(n165, n1417_mux);
buf(g146, n165);
xor (n1418, n1359_mux, n1409_mux);
buf(n1419, n1418_mux);
buf(n166, n1419_mux);
buf(g147, n166);
xor (n1420, n1360_mux, n1408_mux);
buf(n1421, n1420_mux);
buf(n167, n1421_mux);
buf(g148, n167);
xor (n1422, n1361_mux, n1407_mux);
buf(n1423, n1422_mux);
buf(n168, n1423_mux);
buf(g149, n168);
xor (n1424, n1362_mux, n1406_mux);
buf(n1425, n1424_mux);
buf(n169, n1425_mux);
buf(g150, n169);
xor (n1426, n1363_mux, n1405_mux);
buf(n1427, n1426_mux);
buf(n170, n1427_mux);
buf(g151, n170);
xor (n1428, n1348_mux, n1364_mux);
xor (n1429, n1428_mux, n1402_mux);
buf(n1430, n1429_mux);
buf(n171, n1430_mux);
buf(g152, n171);
xor (n1431, n1349_mux, n1365_mux);
xor (n1432, n1431_mux, n1399_mux);
buf(n1433, n1432_mux);
buf(n172, n1433_mux);
buf(g153, n172);
xor (n1434, n1350_mux, n1366_mux);
xor (n1435, n1434_mux, n1396_mux);
buf(n1436, n1435_mux);
buf(n173, n1436_mux);
buf(g154, n173);
xor (n1437, n1351_mux, n1367_mux);
xor (n1438, n1437_mux, n1393_mux);
buf(n1439, n1438_mux);
buf(n174, n1439_mux);
buf(g155, n174);
xor (n1440, n1352_mux, n1368_mux);
xor (n1441, n1440_mux, n1390_mux);
buf(n1442, n1441_mux);
buf(n175, n1442_mux);
buf(g156, n175);
xor (n1443, n1353_mux, n1369_mux);
xor (n1444, n1443_mux, n1387_mux);
buf(n1445, n1444_mux);
buf(n176, n1445_mux);
buf(g157, n176);
xor (n1446, n1354_mux, n1370_mux);
xor (n1447, n1446_mux, n1384_mux);
buf(n1448, n1447_mux);
buf(n177, n1448_mux);
buf(g158, n177);
xor (n1449, n1355_mux, n1371_mux);
xor (n1450, n1449_mux, n1381_mux);
buf(n1451, n1450_mux);
buf(n178, n1451_mux);
buf(g159, n178);
xor (n1452, n1356_mux, n1372_mux);
buf(n1453, n1452_mux);
buf(n179, n1453_mux);
buf(g160, n179);
xor (n852, n654_mux, n657_mux);
xor (n846, n640_mux, n643_mux);
xor (n858, n668_mux, n671_mux);
xor (n861, n675_mux, n678_mux);
xor (n862, n861, n686_mux);
xor (n855, n661_mux, n664_mux);
xor (n856, n855, n692_mux);
xor (n847, n846, n701_mux);
buf(n857, n856);
buf(n848, n847);
xor (n859, n858, n689_mux);
buf(n863, n862);
xor (n853, n852, n695_mux);
xor (n849, n647_mux, n650_mux);
buf(n860, n859);
xor (n864, n682_mux, n685_mux);
buf(n865, n864);
xor (n850, n849, n698_mux);
buf(n851, n850);
buf(n854, n853);
buf(n51, 1'b0);
buf(g32, n51);
buf(n52, 1'b0);
buf(g33, n52);
buf(n53, 1'b0);
buf(g34, n53);
buf(n54, 1'b0);
buf(g35, n54);
buf(n55, 1'b0);
buf(g36, n55);
buf(n56, 1'b0);
buf(g37, n56);
buf(n57, 1'b0);
buf(g38, n57);
buf(n58, 1'b0);
buf(g39, n58);
buf(n59, 1'b0);
buf(g40, n59);
buf(n60, 1'b0);
buf(g41, n60);
buf(n61, 1'b0);
buf(g42, n61);
buf(n62, 1'b0);
buf(g43, n62);
buf(n63, 1'b0);
buf(g44, n63);
buf(n64, 1'b0);
buf(g45, n64);
buf(n65, 1'b0);
buf(g46, n65);
buf(n66, 1'b0);
buf(g47, n66);
buf(n67, 1'b0);
buf(g48, n67);
buf(n68, 1'b0);
buf(g49, n68);
buf(n69, 1'b0);
buf(g50, n69);
buf(n70, 1'b0);
buf(g51, n70);
buf(n71, 1'b0);
buf(g52, n71);
buf(n72, 1'b0);
buf(g53, n72);
buf(n73, 1'b0);
buf(g54, n73);
buf(n74, 1'b0);
buf(g55, n74);
buf(n75, 1'b0);
buf(g56, n75);
buf(n76, 1'b0);
buf(g57, n76);
buf(n77, 1'b0);
buf(g58, n77);
buf(n78, 1'b0);
buf(g59, n78);
buf(n79, 1'b0);
buf(g60, n79);
buf(n80, 1'b0);
buf(g61, n80);
buf(n81, 1'b0);
buf(g62, n81);
buf(n82, 1'b0);
buf(g63, n82);
buf(n83, 1'b0);
buf(g64, n83);
buf(n84, 1'b0);
buf(g65, n84);
buf(n85, 1'b0);
buf(g66, n85);
buf(n86, 1'b0);
buf(g67, n86);
buf(n87, 1'b0);
buf(g68, n87);
buf(n88, 1'b0);
buf(g69, n88);
buf(n89, 1'b0);
buf(g70, n89);
buf(n90, 1'b0);
buf(g71, n90);
buf(n91, 1'b0);
buf(g72, n91);
buf(n92, 1'b0);
buf(g73, n92);
buf(n93, 1'b0);
buf(g74, n93);
buf(n94, 1'b0);
buf(g75, n94);
buf(n95, 1'b0);
buf(g76, n95);
buf(n96, 1'b0);
buf(g77, n96);
buf(n97, 1'b0);
buf(g78, n97);
buf(n98, 1'b0);
buf(g79, n98);
xnor (g0_xnor, g0, g0);
buf(g349, g0_mux);
buf(g349, g0);
xnor (g349_xnor, g349, g349);
buf(n384, g349_mux);
buf(n384, g349);
xnor (n384_xnor, n384, n384);
xnor (g16_xnor, g16, g16);
buf(n35, g16_mux);
buf(n35, g16);
xnor (n35_xnor, n35, n35);
buf(n380, n35_mux);
buf(n380, n35);
xnor (n380_xnor, n380, n380);
and (n1107, n384_mux, n380_mux);
and (n1107, n384, n380);
xnor (n1107_xnor, n1107, n1107);
xnor (g3_xnor, g3, g3);
buf(g352, g3_mux);
buf(g352, g3);
xnor (g352_xnor, g352, g352);
buf(n325, g352_mux);
buf(n325, g352);
xnor (n325_xnor, n325, n325);
not(n1108, n325_mux);
not(n1108, n325);
xnor (n1108_xnor, n1108, n1108);
not(n381, n380_mux);
not(n381, n380);
xnor (n381_xnor, n381, n381);
and (n1109, n381_mux, n325_mux);
and (n1109, n381, n325);
xnor (n1109_xnor, n1109, n1109);
nor (n1110, n1108_mux, n1109_mux);
nor (n1110, n1108, n1109);
xnor (n1110_xnor, n1110, n1110);
xnor (g2_xnor, g2, g2);
buf(g351, g2_mux);
buf(g351, g2);
xnor (g351_xnor, g351, g351);
buf(n334, g351_mux);
buf(n334, g351);
xnor (n334_xnor, n334, n334);
xnor (g17_xnor, g17, g17);
buf(n36, g17_mux);
buf(n36, g17);
xnor (n36_xnor, n36, n36);
buf(n307, n36_mux);
buf(n307, n36);
xnor (n307_xnor, n307, n307);
and (n1111, n334_mux, n307_mux);
and (n1111, n334, n307);
xnor (n1111_xnor, n1111, n1111);
and (n1112, n1110_mux, n1111_mux);
and (n1112, n1110, n1111);
xnor (n1112_xnor, n1112, n1112);
xnor (g1_xnor, g1, g1);
buf(g350, g1_mux);
buf(g350, g1);
xnor (g350_xnor, g350, g350);
buf(n350, g350_mux);
buf(n350, g350);
xnor (n350_xnor, n350, n350);
xnor (g18_xnor, g18, g18);
buf(n37, g18_mux);
buf(n37, g18);
xnor (n37_xnor, n37, n37);
buf(n310, n37_mux);
buf(n310, n37);
xnor (n310_xnor, n310, n310);
and (n1113, n350_mux, n310_mux);
and (n1113, n350, n310);
xnor (n1113_xnor, n1113, n1113);
and (n1114, n1111_mux, n1113_mux);
and (n1114, n1111, n1113);
xnor (n1114_xnor, n1114, n1114);
and (n1115, n1110_mux, n1113_mux);
and (n1115, n1110, n1113);
xnor (n1115_xnor, n1115, n1115);
or (n1116_1, n1114_mux, n1115_mux);
or (n1116, n1112_mux, n1116_1);
or (n1116_1, n1114, n1115);
or (n1116, n1112, n1116_1);
xnor (n1116_xnor, n1116, n1116);
not(n1117, n334_mux);
not(n1117, n334);
xnor (n1117_xnor, n1117, n1117);
and (n1118, n381_mux, n334_mux);
and (n1118, n381, n334);
xnor (n1118_xnor, n1118, n1118);
nor (n1119, n1117_mux, n1118_mux);
nor (n1119, n1117, n1118);
xnor (n1119_xnor, n1119, n1119);
and (n1120, n1116_mux, n1119_mux);
and (n1120, n1116, n1119);
xnor (n1120_xnor, n1120, n1120);
and (n1121, n350_mux, n307_mux);
and (n1121, n350, n307);
xnor (n1121_xnor, n1121, n1121);
and (n1122, n1119_mux, n1121_mux);
and (n1122, n1119, n1121);
xnor (n1122_xnor, n1122, n1122);
and (n1123, n1116_mux, n1121_mux);
and (n1123, n1116, n1121);
xnor (n1123_xnor, n1123, n1123);
or (n1124_1, n1122_mux, n1123_mux);
or (n1124, n1120_mux, n1124_1);
or (n1124_1, n1122, n1123);
or (n1124, n1120, n1124_1);
xnor (n1124_xnor, n1124, n1124);
not(n1125, n350_mux);
not(n1125, n350);
xnor (n1125_xnor, n1125, n1125);
and (n1126, n381_mux, n350_mux);
and (n1126, n381, n350);
xnor (n1126_xnor, n1126, n1126);
nor (n1127, n1125_mux, n1126_mux);
nor (n1127, n1125, n1126);
xnor (n1127_xnor, n1127, n1127);
and (n1128, n1124_mux, n1127_mux);
and (n1128, n1124, n1127);
xnor (n1128_xnor, n1128, n1128);
not(n385, n384_mux);
not(n385, n384);
xnor (n385_xnor, n385, n385);
and (n1129, n385_mux, n307_mux);
and (n1129, n385, n307);
xnor (n1129_xnor, n1129, n1129);
not(n1130, n307_mux);
not(n1130, n307);
xnor (n1130_xnor, n1130, n1130);
nor (n1131, n1129_mux, n1130_mux);
nor (n1131, n1129, n1130);
xnor (n1131_xnor, n1131, n1131);
and (n1132, n1127_mux, n1131_mux);
and (n1132, n1127, n1131);
xnor (n1132_xnor, n1132, n1132);
and (n1133, n1124_mux, n1131_mux);
and (n1133, n1124, n1131);
xnor (n1133_xnor, n1133, n1133);
or (n1134_1, n1132_mux, n1133_mux);
or (n1134, n1128_mux, n1134_1);
or (n1134_1, n1132, n1133);
or (n1134, n1128, n1134_1);
xnor (n1134_xnor, n1134, n1134);
and (n1135, n1107_mux, n1134_mux);
and (n1135, n1107, n1134);
xnor (n1135_xnor, n1135, n1135);
xor (n1136, n1107_mux, n1134_mux);
xor (n1136, n1107, n1134);
xnor (n1136_xnor, n1136, n1136);
xor (n1137, n1124_mux, n1127_mux);
xor (n1137, n1124, n1127);
xnor (n1137_xnor, n1137, n1137);
xor (n1138, n1137_mux, n1131_mux);
xor (n1138, n1137, n1131);
xnor (n1138_xnor, n1138, n1138);
xnor (g4_xnor, g4, g4);
buf(g353, g4_mux);
buf(g353, g4);
xnor (g353_xnor, g353, g353);
buf(n321, g353_mux);
buf(n321, g353);
xnor (n321_xnor, n321, n321);
not(n1139, n321_mux);
not(n1139, n321);
xnor (n1139_xnor, n1139, n1139);
and (n1140, n381_mux, n321_mux);
and (n1140, n381, n321);
xnor (n1140_xnor, n1140, n1140);
nor (n1141, n1139_mux, n1140_mux);
nor (n1141, n1139, n1140);
xnor (n1141_xnor, n1141, n1141);
and (n1142, n325_mux, n307_mux);
and (n1142, n325, n307);
xnor (n1142_xnor, n1142, n1142);
and (n1143, n1141_mux, n1142_mux);
and (n1143, n1141, n1142);
xnor (n1143_xnor, n1143, n1143);
xnor (g20_xnor, g20, g20);
buf(n39, g20_mux);
buf(n39, g20);
xnor (n39_xnor, n39, n39);
buf(n344, n39_mux);
buf(n344, n39);
xnor (n344_xnor, n344, n344);
and (n1144, n385_mux, n344_mux);
and (n1144, n385, n344);
xnor (n1144_xnor, n1144, n1144);
not(n1145, n344_mux);
not(n1145, n344);
xnor (n1145_xnor, n1145, n1145);
nor (n1146, n1144_mux, n1145_mux);
nor (n1146, n1144, n1145);
xnor (n1146_xnor, n1146, n1146);
and (n1147, n1142_mux, n1146_mux);
and (n1147, n1142, n1146);
xnor (n1147_xnor, n1147, n1147);
and (n1148, n1141_mux, n1146_mux);
and (n1148, n1141, n1146);
xnor (n1148_xnor, n1148, n1148);
or (n1149_1, n1147_mux, n1148_mux);
or (n1149, n1143_mux, n1149_1);
or (n1149_1, n1147, n1148);
or (n1149, n1143, n1149_1);
xnor (n1149_xnor, n1149, n1149);
and (n1150, n325_mux, n310_mux);
and (n1150, n325, n310);
xnor (n1150_xnor, n1150, n1150);
xnor (g19_xnor, g19, g19);
buf(n38, g19_mux);
buf(n38, g19);
xnor (n38_xnor, n38, n38);
buf(n314, n38_mux);
buf(n314, n38);
xnor (n314_xnor, n314, n314);
and (n1151, n334_mux, n314_mux);
and (n1151, n334, n314);
xnor (n1151_xnor, n1151, n1151);
and (n1152, n1150_mux, n1151_mux);
and (n1152, n1150, n1151);
xnor (n1152_xnor, n1152, n1152);
and (n1153, n350_mux, n344_mux);
and (n1153, n350, n344);
xnor (n1153_xnor, n1153, n1153);
and (n1154, n1151_mux, n1153_mux);
and (n1154, n1151, n1153);
xnor (n1154_xnor, n1154, n1154);
and (n1155, n1150_mux, n1153_mux);
and (n1155, n1150, n1153);
xnor (n1155_xnor, n1155, n1155);
or (n1156_1, n1154_mux, n1155_mux);
or (n1156, n1152_mux, n1156_1);
or (n1156_1, n1154, n1155);
or (n1156, n1152, n1156_1);
xnor (n1156_xnor, n1156, n1156);
and (n1157, n334_mux, n310_mux);
and (n1157, n334, n310);
xnor (n1157_xnor, n1157, n1157);
and (n1158, n1156_mux, n1157_mux);
and (n1158, n1156, n1157);
xnor (n1158_xnor, n1158, n1158);
and (n1159, n350_mux, n314_mux);
and (n1159, n350, n314);
xnor (n1159_xnor, n1159, n1159);
and (n1160, n1157_mux, n1159_mux);
and (n1160, n1157, n1159);
xnor (n1160_xnor, n1160, n1160);
and (n1161, n1156_mux, n1159_mux);
and (n1161, n1156, n1159);
xnor (n1161_xnor, n1161, n1161);
or (n1162_1, n1160_mux, n1161_mux);
or (n1162, n1158_mux, n1162_1);
or (n1162_1, n1160, n1161);
or (n1162, n1158, n1162_1);
xnor (n1162_xnor, n1162, n1162);
and (n1163, n1149_mux, n1162_mux);
and (n1163, n1149, n1162);
xnor (n1163_xnor, n1163, n1163);
xor (n1164, n1110_mux, n1111_mux);
xor (n1164, n1110, n1111);
xnor (n1164_xnor, n1164, n1164);
xor (n1165, n1164_mux, n1113_mux);
xor (n1165, n1164, n1113);
xnor (n1165_xnor, n1165, n1165);
and (n1166, n1162_mux, n1165_mux);
and (n1166, n1162, n1165);
xnor (n1166_xnor, n1166, n1166);
and (n1167, n1149_mux, n1165_mux);
and (n1167, n1149, n1165);
xnor (n1167_xnor, n1167, n1167);
or (n1168_1, n1166_mux, n1167_mux);
or (n1168, n1163_mux, n1168_1);
or (n1168_1, n1166, n1167);
or (n1168, n1163, n1168_1);
xnor (n1168_xnor, n1168, n1168);
and (n1169, n385_mux, n310_mux);
and (n1169, n385, n310);
xnor (n1169_xnor, n1169, n1169);
not(n1170, n310_mux);
not(n1170, n310);
xnor (n1170_xnor, n1170, n1170);
nor (n1171, n1169_mux, n1170_mux);
nor (n1171, n1169, n1170);
xnor (n1171_xnor, n1171, n1171);
and (n1172, n1168_mux, n1171_mux);
and (n1172, n1168, n1171);
xnor (n1172_xnor, n1172, n1172);
xor (n1173, n1116_mux, n1119_mux);
xor (n1173, n1116, n1119);
xnor (n1173_xnor, n1173, n1173);
xor (n1174, n1173_mux, n1121_mux);
xor (n1174, n1173, n1121);
xnor (n1174_xnor, n1174, n1174);
and (n1175, n1171_mux, n1174_mux);
and (n1175, n1171, n1174);
xnor (n1175_xnor, n1175, n1175);
and (n1176, n1168_mux, n1174_mux);
and (n1176, n1168, n1174);
xnor (n1176_xnor, n1176, n1176);
or (n1177_1, n1175_mux, n1176_mux);
or (n1177, n1172_mux, n1177_1);
or (n1177_1, n1175, n1176);
or (n1177, n1172, n1177_1);
xnor (n1177_xnor, n1177, n1177);
and (n1178, n1138_mux, n1177_mux);
and (n1178, n1138, n1177);
xnor (n1178_xnor, n1178, n1178);
xor (n1179, n1138_mux, n1177_mux);
xor (n1179, n1138, n1177);
xnor (n1179_xnor, n1179, n1179);
xor (n1180, n1168_mux, n1171_mux);
xor (n1180, n1168, n1171);
xnor (n1180_xnor, n1180, n1180);
xor (n1181, n1180_mux, n1174_mux);
xor (n1181, n1180, n1174);
xnor (n1181_xnor, n1181, n1181);
and (n1182, n325_mux, n314_mux);
and (n1182, n325, n314);
xnor (n1182_xnor, n1182, n1182);
and (n1183, n334_mux, n344_mux);
and (n1183, n334, n344);
xnor (n1183_xnor, n1183, n1183);
and (n1184, n1182_mux, n1183_mux);
and (n1184, n1182, n1183);
xnor (n1184_xnor, n1184, n1184);
xnor (g21_xnor, g21, g21);
buf(n40, g21_mux);
buf(n40, g21);
xnor (n40_xnor, n40, n40);
buf(n319, n40_mux);
buf(n319, n40);
xnor (n319_xnor, n319, n319);
and (n1185, n350_mux, n319_mux);
and (n1185, n350, n319);
xnor (n1185_xnor, n1185, n1185);
and (n1186, n1183_mux, n1185_mux);
and (n1186, n1183, n1185);
xnor (n1186_xnor, n1186, n1186);
and (n1187, n1182_mux, n1185_mux);
and (n1187, n1182, n1185);
xnor (n1187_xnor, n1187, n1187);
or (n1188_1, n1186_mux, n1187_mux);
or (n1188, n1184_mux, n1188_1);
or (n1188_1, n1186, n1187);
or (n1188, n1184, n1188_1);
xnor (n1188_xnor, n1188, n1188);
xnor (g5_xnor, g5, g5);
buf(g354, g5_mux);
buf(g354, g5);
xnor (g354_xnor, g354, g354);
buf(n313, g354_mux);
buf(n313, g354);
xnor (n313_xnor, n313, n313);
and (n1189, n313_mux, n307_mux);
and (n1189, n313, n307);
xnor (n1189_xnor, n1189, n1189);
and (n1190, n321_mux, n310_mux);
and (n1190, n321, n310);
xnor (n1190_xnor, n1190, n1190);
and (n1191, n1189_mux, n1190_mux);
and (n1191, n1189, n1190);
xnor (n1191_xnor, n1191, n1191);
and (n1192, n1188_mux, n1191_mux);
and (n1192, n1188, n1191);
xnor (n1192_xnor, n1192, n1192);
xor (n1193, n1150_mux, n1151_mux);
xor (n1193, n1150, n1151);
xnor (n1193_xnor, n1193, n1193);
xor (n1194, n1193_mux, n1153_mux);
xor (n1194, n1193, n1153);
xnor (n1194_xnor, n1194, n1194);
and (n1195, n1191_mux, n1194_mux);
and (n1195, n1191, n1194);
xnor (n1195_xnor, n1195, n1195);
and (n1196, n1188_mux, n1194_mux);
and (n1196, n1188, n1194);
xnor (n1196_xnor, n1196, n1196);
or (n1197_1, n1195_mux, n1196_mux);
or (n1197, n1192_mux, n1197_1);
or (n1197_1, n1195, n1196);
or (n1197, n1192, n1197_1);
xnor (n1197_xnor, n1197, n1197);
xor (n1198, n1141_mux, n1142_mux);
xor (n1198, n1141, n1142);
xnor (n1198_xnor, n1198, n1198);
xor (n1199, n1198_mux, n1146_mux);
xor (n1199, n1198, n1146);
xnor (n1199_xnor, n1199, n1199);
and (n1200, n1197_mux, n1199_mux);
and (n1200, n1197, n1199);
xnor (n1200_xnor, n1200, n1200);
xor (n1201, n1156_mux, n1157_mux);
xor (n1201, n1156, n1157);
xnor (n1201_xnor, n1201, n1201);
xor (n1202, n1201_mux, n1159_mux);
xor (n1202, n1201, n1159);
xnor (n1202_xnor, n1202, n1202);
and (n1203, n1199_mux, n1202_mux);
and (n1203, n1199, n1202);
xnor (n1203_xnor, n1203, n1203);
and (n1204, n1197_mux, n1202_mux);
and (n1204, n1197, n1202);
xnor (n1204_xnor, n1204, n1204);
or (n1205_1, n1203_mux, n1204_mux);
or (n1205, n1200_mux, n1205_1);
or (n1205_1, n1203, n1204);
or (n1205, n1200, n1205_1);
xnor (n1205_xnor, n1205, n1205);
and (n1206, n385_mux, n314_mux);
and (n1206, n385, n314);
xnor (n1206_xnor, n1206, n1206);
not(n1207, n314_mux);
not(n1207, n314);
xnor (n1207_xnor, n1207, n1207);
nor (n1208, n1206_mux, n1207_mux);
nor (n1208, n1206, n1207);
xnor (n1208_xnor, n1208, n1208);
and (n1209, n1205_mux, n1208_mux);
and (n1209, n1205, n1208);
xnor (n1209_xnor, n1209, n1209);
xor (n1210, n1149_mux, n1162_mux);
xor (n1210, n1149, n1162);
xnor (n1210_xnor, n1210, n1210);
xor (n1211, n1210_mux, n1165_mux);
xor (n1211, n1210, n1165);
xnor (n1211_xnor, n1211, n1211);
and (n1212, n1208_mux, n1211_mux);
and (n1212, n1208, n1211);
xnor (n1212_xnor, n1212, n1212);
and (n1213, n1205_mux, n1211_mux);
and (n1213, n1205, n1211);
xnor (n1213_xnor, n1213, n1213);
or (n1214_1, n1212_mux, n1213_mux);
or (n1214, n1209_mux, n1214_1);
or (n1214_1, n1212, n1213);
or (n1214, n1209, n1214_1);
xnor (n1214_xnor, n1214, n1214);
and (n1215, n1181_mux, n1214_mux);
and (n1215, n1181, n1214);
xnor (n1215_xnor, n1215, n1215);
xor (n1216, n1181_mux, n1214_mux);
xor (n1216, n1181, n1214);
xnor (n1216_xnor, n1216, n1216);
xor (n1217, n1205_mux, n1208_mux);
xor (n1217, n1205, n1208);
xnor (n1217_xnor, n1217, n1217);
xor (n1218, n1217_mux, n1211_mux);
xor (n1218, n1217, n1211);
xnor (n1218_xnor, n1218, n1218);
not(n1219, n313_mux);
not(n1219, n313);
xnor (n1219_xnor, n1219, n1219);
and (n1220, n381_mux, n313_mux);
and (n1220, n381, n313);
xnor (n1220_xnor, n1220, n1220);
nor (n1221, n1219_mux, n1220_mux);
nor (n1221, n1219, n1220);
xnor (n1221_xnor, n1221, n1221);
and (n1222, n321_mux, n307_mux);
and (n1222, n321, n307);
xnor (n1222_xnor, n1222, n1222);
and (n1223, n1221_mux, n1222_mux);
and (n1223, n1221, n1222);
xnor (n1223_xnor, n1223, n1223);
and (n1224, n385_mux, n319_mux);
and (n1224, n385, n319);
xnor (n1224_xnor, n1224, n1224);
not(n1225, n319_mux);
not(n1225, n319);
xnor (n1225_xnor, n1225, n1225);
nor (n1226, n1224_mux, n1225_mux);
nor (n1226, n1224, n1225);
xnor (n1226_xnor, n1226, n1226);
and (n1227, n1222_mux, n1226_mux);
and (n1227, n1222, n1226);
xnor (n1227_xnor, n1227, n1227);
and (n1228, n1221_mux, n1226_mux);
and (n1228, n1221, n1226);
xnor (n1228_xnor, n1228, n1228);
or (n1229_1, n1227_mux, n1228_mux);
or (n1229, n1223_mux, n1229_1);
or (n1229_1, n1227, n1228);
or (n1229, n1223, n1229_1);
xnor (n1229_xnor, n1229, n1229);
and (n372, n325_mux, n344_mux);
and (n372, n325, n344);
xnor (n372_xnor, n372, n372);
and (n373, n334_mux, n319_mux);
and (n373, n334, n319);
xnor (n373_xnor, n373, n373);
and (n1230, n372_mux, n373_mux);
and (n1230, n372, n373);
xnor (n1230_xnor, n1230, n1230);
xnor (g22_xnor, g22, g22);
buf(n41, g22_mux);
buf(n41, g22);
xnor (n41_xnor, n41, n41);
buf(n322, n41_mux);
buf(n322, n41);
xnor (n322_xnor, n322, n322);
and (n375, n350_mux, n322_mux);
and (n375, n350, n322);
xnor (n375_xnor, n375, n375);
and (n1231, n373_mux, n375_mux);
and (n1231, n373, n375);
xnor (n1231_xnor, n1231, n1231);
and (n1232, n372_mux, n375_mux);
and (n1232, n372, n375);
xnor (n1232_xnor, n1232, n1232);
or (n1233_1, n1231_mux, n1232_mux);
or (n1233, n1230_mux, n1233_1);
or (n1233_1, n1231, n1232);
or (n1233, n1230, n1233_1);
xnor (n1233_xnor, n1233, n1233);
xor (n1234, n1182_mux, n1183_mux);
xor (n1234, n1182, n1183);
xnor (n1234_xnor, n1234, n1234);
xor (n1235, n1234_mux, n1185_mux);
xor (n1235, n1234, n1185);
xnor (n1235_xnor, n1235, n1235);
and (n1236, n1233_mux, n1235_mux);
and (n1236, n1233, n1235);
xnor (n1236_xnor, n1236, n1236);
xor (n1237, n1189_mux, n1190_mux);
xor (n1237, n1189, n1190);
xnor (n1237_xnor, n1237, n1237);
and (n1238, n1235_mux, n1237_mux);
and (n1238, n1235, n1237);
xnor (n1238_xnor, n1238, n1238);
and (n1239, n1233_mux, n1237_mux);
and (n1239, n1233, n1237);
xnor (n1239_xnor, n1239, n1239);
or (n1240_1, n1238_mux, n1239_mux);
or (n1240, n1236_mux, n1240_1);
or (n1240_1, n1238, n1239);
or (n1240, n1236, n1240_1);
xnor (n1240_xnor, n1240, n1240);
xor (n1241, n1221_mux, n1222_mux);
xor (n1241, n1221, n1222);
xnor (n1241_xnor, n1241, n1241);
xor (n1242, n1241_mux, n1226_mux);
xor (n1242, n1241, n1226);
xnor (n1242_xnor, n1242, n1242);
and (n1243, n1240_mux, n1242_mux);
and (n1243, n1240, n1242);
xnor (n1243_xnor, n1243, n1243);
xor (n1244, n1188_mux, n1191_mux);
xor (n1244, n1188, n1191);
xnor (n1244_xnor, n1244, n1244);
xor (n1245, n1244_mux, n1194_mux);
xor (n1245, n1244, n1194);
xnor (n1245_xnor, n1245, n1245);
and (n1246, n1242_mux, n1245_mux);
and (n1246, n1242, n1245);
xnor (n1246_xnor, n1246, n1246);
and (n1247, n1240_mux, n1245_mux);
and (n1247, n1240, n1245);
xnor (n1247_xnor, n1247, n1247);
or (n1248_1, n1246_mux, n1247_mux);
or (n1248, n1243_mux, n1248_1);
or (n1248_1, n1246, n1247);
or (n1248, n1243, n1248_1);
xnor (n1248_xnor, n1248, n1248);
and (n1249, n1229_mux, n1248_mux);
and (n1249, n1229, n1248);
xnor (n1249_xnor, n1249, n1249);
xor (n1250, n1197_mux, n1199_mux);
xor (n1250, n1197, n1199);
xnor (n1250_xnor, n1250, n1250);
xor (n1251, n1250_mux, n1202_mux);
xor (n1251, n1250, n1202);
xnor (n1251_xnor, n1251, n1251);
and (n1252, n1248_mux, n1251_mux);
and (n1252, n1248, n1251);
xnor (n1252_xnor, n1252, n1252);
and (n1253, n1229_mux, n1251_mux);
and (n1253, n1229, n1251);
xnor (n1253_xnor, n1253, n1253);
or (n1254_1, n1252_mux, n1253_mux);
or (n1254, n1249_mux, n1254_1);
or (n1254_1, n1252, n1253);
or (n1254, n1249, n1254_1);
xnor (n1254_xnor, n1254, n1254);
and (n1255, n1218_mux, n1254_mux);
and (n1255, n1218, n1254);
xnor (n1255_xnor, n1255, n1255);
xor (n1256, n1218_mux, n1254_mux);
xor (n1256, n1218, n1254);
xnor (n1256_xnor, n1256, n1256);
xor (n1257, n1229_mux, n1248_mux);
xor (n1257, n1229, n1248);
xnor (n1257_xnor, n1257, n1257);
xor (n1258, n1257_mux, n1251_mux);
xor (n1258, n1257, n1251);
xnor (n1258_xnor, n1258, n1258);
xnor (g6_xnor, g6, g6);
buf(g355, g6_mux);
buf(g355, g6);
xnor (g355_xnor, g355, g355);
buf(n309, g355_mux);
buf(n309, g355);
xnor (n309_xnor, n309, n309);
and (n366, n309_mux, n307_mux);
and (n366, n309, n307);
xnor (n366_xnor, n366, n366);
and (n367, n313_mux, n310_mux);
and (n367, n313, n310);
xnor (n367_xnor, n367, n367);
and (n1259, n366_mux, n367_mux);
and (n1259, n366, n367);
xnor (n1259_xnor, n1259, n1259);
and (n369, n321_mux, n314_mux);
and (n369, n321, n314);
xnor (n369_xnor, n369, n369);
and (n1260, n367_mux, n369_mux);
and (n1260, n367, n369);
xnor (n1260_xnor, n1260, n1260);
and (n1261, n366_mux, n369_mux);
and (n1261, n366, n369);
xnor (n1261_xnor, n1261, n1261);
or (n1262_1, n1260_mux, n1261_mux);
or (n1262, n1259_mux, n1262_1);
or (n1262_1, n1260, n1261);
or (n1262, n1259, n1262_1);
xnor (n1262_xnor, n1262, n1262);
not(n1263, n309_mux);
not(n1263, n309);
xnor (n1263_xnor, n1263, n1263);
and (n1264, n381_mux, n309_mux);
and (n1264, n381, n309);
xnor (n1264_xnor, n1264, n1264);
nor (n1265, n1263_mux, n1264_mux);
nor (n1265, n1263, n1264);
xnor (n1265_xnor, n1265, n1265);
and (n1266, n1262_mux, n1265_mux);
and (n1266, n1262, n1265);
xnor (n1266_xnor, n1266, n1266);
and (n1267, n385_mux, n322_mux);
and (n1267, n385, n322);
xnor (n1267_xnor, n1267, n1267);
not(n1268, n322_mux);
not(n1268, n322);
xnor (n1268_xnor, n1268, n1268);
nor (n1269, n1267_mux, n1268_mux);
nor (n1269, n1267, n1268);
xnor (n1269_xnor, n1269, n1269);
and (n1270, n1265_mux, n1269_mux);
and (n1270, n1265, n1269);
xnor (n1270_xnor, n1270, n1270);
and (n1271, n1262_mux, n1269_mux);
and (n1271, n1262, n1269);
xnor (n1271_xnor, n1271, n1271);
or (n1272_1, n1270_mux, n1271_mux);
or (n1272, n1266_mux, n1272_1);
or (n1272_1, n1270, n1271);
or (n1272, n1266, n1272_1);
xnor (n1272_xnor, n1272, n1272);
and (n347, n325_mux, n319_mux);
and (n347, n325, n319);
xnor (n347_xnor, n347, n347);
and (n348, n334_mux, n322_mux);
and (n348, n334, n322);
xnor (n348_xnor, n348, n348);
and (n362, n347_mux, n348_mux);
and (n362, n347, n348);
xnor (n362_xnor, n362, n362);
xnor (g23_xnor, g23, g23);
buf(n42, g23_mux);
buf(n42, g23);
xnor (n42_xnor, n42, n42);
buf(n326, n42_mux);
buf(n326, n42);
xnor (n326_xnor, n326, n326);
and (n351, n350_mux, n326_mux);
and (n351, n350, n326);
xnor (n351_xnor, n351, n351);
and (n363, n348_mux, n351_mux);
and (n363, n348, n351);
xnor (n363_xnor, n363, n363);
and (n364, n347_mux, n351_mux);
and (n364, n347, n351);
xnor (n364_xnor, n364, n364);
or (n365_1, n363_mux, n364_mux);
or (n365, n362_mux, n365_1);
or (n365_1, n363, n364);
or (n365, n362, n365_1);
xnor (n365_xnor, n365, n365);
xor (n368, n366_mux, n367_mux);
xor (n368, n366, n367);
xnor (n368_xnor, n368, n368);
xor (n370, n368_mux, n369_mux);
xor (n370, n368, n369);
xnor (n370_xnor, n370, n370);
and (n1273, n365_mux, n370_mux);
and (n1273, n365, n370);
xnor (n1273_xnor, n1273, n1273);
xor (n374, n372_mux, n373_mux);
xor (n374, n372, n373);
xnor (n374_xnor, n374, n374);
xor (n376, n374_mux, n375_mux);
xor (n376, n374, n375);
xnor (n376_xnor, n376, n376);
and (n1274, n370_mux, n376_mux);
and (n1274, n370, n376);
xnor (n1274_xnor, n1274, n1274);
and (n1275, n365_mux, n376_mux);
and (n1275, n365, n376);
xnor (n1275_xnor, n1275, n1275);
or (n1276_1, n1274_mux, n1275_mux);
or (n1276, n1273_mux, n1276_1);
or (n1276_1, n1274, n1275);
or (n1276, n1273, n1276_1);
xnor (n1276_xnor, n1276, n1276);
xor (n1277, n1262_mux, n1265_mux);
xor (n1277, n1262, n1265);
xnor (n1277_xnor, n1277, n1277);
xor (n1278, n1277_mux, n1269_mux);
xor (n1278, n1277, n1269);
xnor (n1278_xnor, n1278, n1278);
and (n1279, n1276_mux, n1278_mux);
and (n1279, n1276, n1278);
xnor (n1279_xnor, n1279, n1279);
xor (n1280, n1233_mux, n1235_mux);
xor (n1280, n1233, n1235);
xnor (n1280_xnor, n1280, n1280);
xor (n1281, n1280_mux, n1237_mux);
xor (n1281, n1280, n1237);
xnor (n1281_xnor, n1281, n1281);
and (n1282, n1278_mux, n1281_mux);
and (n1282, n1278, n1281);
xnor (n1282_xnor, n1282, n1282);
and (n1283, n1276_mux, n1281_mux);
and (n1283, n1276, n1281);
xnor (n1283_xnor, n1283, n1283);
or (n1284_1, n1282_mux, n1283_mux);
or (n1284, n1279_mux, n1284_1);
or (n1284_1, n1282, n1283);
or (n1284, n1279, n1284_1);
xnor (n1284_xnor, n1284, n1284);
and (n1285, n1272_mux, n1284_mux);
and (n1285, n1272, n1284);
xnor (n1285_xnor, n1285, n1285);
xor (n1286, n1240_mux, n1242_mux);
xor (n1286, n1240, n1242);
xnor (n1286_xnor, n1286, n1286);
xor (n1287, n1286_mux, n1245_mux);
xor (n1287, n1286, n1245);
xnor (n1287_xnor, n1287, n1287);
and (n1288, n1284_mux, n1287_mux);
and (n1288, n1284, n1287);
xnor (n1288_xnor, n1288, n1288);
and (n1289, n1272_mux, n1287_mux);
and (n1289, n1272, n1287);
xnor (n1289_xnor, n1289, n1289);
or (n1290_1, n1288_mux, n1289_mux);
or (n1290, n1285_mux, n1290_1);
or (n1290_1, n1288, n1289);
or (n1290, n1285, n1290_1);
xnor (n1290_xnor, n1290, n1290);
and (n1291, n1258_mux, n1290_mux);
and (n1291, n1258, n1290);
xnor (n1291_xnor, n1291, n1291);
xor (n1292, n1258_mux, n1290_mux);
xor (n1292, n1258, n1290);
xnor (n1292_xnor, n1292, n1292);
xor (n1293, n1272_mux, n1284_mux);
xor (n1293, n1272, n1284);
xnor (n1293_xnor, n1293, n1293);
xor (n1294, n1293_mux, n1287_mux);
xor (n1294, n1293, n1287);
xnor (n1294_xnor, n1294, n1294);
xnor (g7_xnor, g7, g7);
buf(g356, g7_mux);
buf(g356, g7);
xnor (g356_xnor, g356, g356);
buf(n306, g356_mux);
buf(n306, g356);
xnor (n306_xnor, n306, n306);
not(n379, n306_mux);
not(n379, n306);
xnor (n379_xnor, n379, n379);
and (n382, n381_mux, n306_mux);
and (n382, n381, n306);
xnor (n382_xnor, n382, n382);
nor (n383, n379_mux, n382_mux);
nor (n383, n379, n382);
xnor (n383_xnor, n383, n383);
and (n386, n385_mux, n326_mux);
and (n386, n385, n326);
xnor (n386_xnor, n386, n386);
not(n387, n326_mux);
not(n387, n326);
xnor (n387_xnor, n387, n387);
nor (n388, n386_mux, n387_mux);
nor (n388, n386, n387);
xnor (n388_xnor, n388, n388);
and (n1295, n383_mux, n388_mux);
and (n1295, n383, n388);
xnor (n1295_xnor, n1295, n1295);
and (n333, n325_mux, n322_mux);
and (n333, n325, n322);
xnor (n333_xnor, n333, n333);
and (n335, n334_mux, n326_mux);
and (n335, n334, n326);
xnor (n335_xnor, n335, n335);
and (n343, n333_mux, n335_mux);
and (n343, n333, n335);
xnor (n343_xnor, n343, n343);
and (n345, n321_mux, n344_mux);
and (n345, n321, n344);
xnor (n345_xnor, n345, n345);
and (n358, n343_mux, n345_mux);
and (n358, n343, n345);
xnor (n358_xnor, n358, n358);
xor (n349, n347_mux, n348_mux);
xor (n349, n347, n348);
xnor (n349_xnor, n349, n349);
xor (n352, n349_mux, n351_mux);
xor (n352, n349, n351);
xnor (n352_xnor, n352, n352);
and (n359, n345_mux, n352_mux);
and (n359, n345, n352);
xnor (n359_xnor, n359, n359);
and (n360, n343_mux, n352_mux);
and (n360, n343, n352);
xnor (n360_xnor, n360, n360);
or (n361_1, n359_mux, n360_mux);
or (n361, n358_mux, n361_1);
or (n361_1, n359, n360);
or (n361, n358, n361_1);
xnor (n361_xnor, n361, n361);
xor (n371, n365_mux, n370_mux);
xor (n371, n365, n370);
xnor (n371_xnor, n371, n371);
xor (n377, n371_mux, n376_mux);
xor (n377, n371, n376);
xnor (n377_xnor, n377, n377);
and (n1296, n361_mux, n377_mux);
and (n1296, n361, n377);
xnor (n1296_xnor, n1296, n1296);
xor (n389, n383_mux, n388_mux);
xor (n389, n383, n388);
xnor (n389_xnor, n389, n389);
and (n1297, n377_mux, n389_mux);
and (n1297, n377, n389);
xnor (n1297_xnor, n1297, n1297);
and (n1298, n361_mux, n389_mux);
and (n1298, n361, n389);
xnor (n1298_xnor, n1298, n1298);
or (n1299_1, n1297_mux, n1298_mux);
or (n1299, n1296_mux, n1299_1);
or (n1299_1, n1297, n1298);
or (n1299, n1296, n1299_1);
xnor (n1299_xnor, n1299, n1299);
and (n1300, n1295_mux, n1299_mux);
and (n1300, n1295, n1299);
xnor (n1300_xnor, n1300, n1300);
xor (n1301, n1276_mux, n1278_mux);
xor (n1301, n1276, n1278);
xnor (n1301_xnor, n1301, n1301);
xor (n1302, n1301_mux, n1281_mux);
xor (n1302, n1301, n1281);
xnor (n1302_xnor, n1302, n1302);
and (n1303, n1299_mux, n1302_mux);
and (n1303, n1299, n1302);
xnor (n1303_xnor, n1303, n1303);
and (n1304, n1295_mux, n1302_mux);
and (n1304, n1295, n1302);
xnor (n1304_xnor, n1304, n1304);
or (n1305_1, n1303_mux, n1304_mux);
or (n1305, n1300_mux, n1305_1);
or (n1305_1, n1303, n1304);
or (n1305, n1300, n1305_1);
xnor (n1305_xnor, n1305, n1305);
and (n1306, n1294_mux, n1305_mux);
and (n1306, n1294, n1305);
xnor (n1306_xnor, n1306, n1306);
xor (n1307, n1294_mux, n1305_mux);
xor (n1307, n1294, n1305);
xnor (n1307_xnor, n1307, n1307);
xor (n1308, n1295_mux, n1299_mux);
xor (n1308, n1295, n1299);
xnor (n1308_xnor, n1308, n1308);
xor (n1309, n1308_mux, n1302_mux);
xor (n1309, n1308, n1302);
xnor (n1309_xnor, n1309, n1309);
and (n308, n306_mux, n307_mux);
and (n308, n306, n307);
xnor (n308_xnor, n308, n308);
and (n311, n309_mux, n310_mux);
and (n311, n309, n310);
xnor (n311_xnor, n311, n311);
and (n312, n308_mux, n311_mux);
and (n312, n308, n311);
xnor (n312_xnor, n312, n312);
and (n315, n313_mux, n314_mux);
and (n315, n313, n314);
xnor (n315_xnor, n315, n315);
and (n316, n311_mux, n315_mux);
and (n316, n311, n315);
xnor (n316_xnor, n316, n316);
and (n317, n308_mux, n315_mux);
and (n317, n308, n315);
xnor (n317_xnor, n317, n317);
or (n318_1, n316_mux, n317_mux);
or (n318, n312_mux, n318_1);
or (n318_1, n316, n317);
or (n318, n312, n318_1);
xnor (n318_xnor, n318, n318);
and (n320, n313_mux, n319_mux);
and (n320, n313, n319);
xnor (n320_xnor, n320, n320);
and (n323, n321_mux, n322_mux);
and (n323, n321, n322);
xnor (n323_xnor, n323, n323);
and (n324, n320_mux, n323_mux);
and (n324, n320, n323);
xnor (n324_xnor, n324, n324);
and (n327, n325_mux, n326_mux);
and (n327, n325, n326);
xnor (n327_xnor, n327, n327);
and (n328, n323_mux, n327_mux);
and (n328, n323, n327);
xnor (n328_xnor, n328, n328);
and (n329, n320_mux, n327_mux);
and (n329, n320, n327);
xnor (n329_xnor, n329, n329);
or (n330_1, n328_mux, n329_mux);
or (n330, n324_mux, n330_1);
or (n330_1, n328, n329);
or (n330, n324, n330_1);
xnor (n330_xnor, n330, n330);
and (n331, n321_mux, n319_mux);
and (n331, n321, n319);
xnor (n331_xnor, n331, n331);
and (n332, n330_mux, n331_mux);
and (n332, n330, n331);
xnor (n332_xnor, n332, n332);
xor (n336, n333_mux, n335_mux);
xor (n336, n333, n335);
xnor (n336_xnor, n336, n336);
and (n337, n331_mux, n336_mux);
and (n337, n331, n336);
xnor (n337_xnor, n337, n337);
and (n338, n330_mux, n336_mux);
and (n338, n330, n336);
xnor (n338_xnor, n338, n338);
or (n339_1, n337_mux, n338_mux);
or (n339, n332_mux, n339_1);
or (n339_1, n337, n338);
or (n339, n332, n339_1);
xnor (n339_xnor, n339, n339);
xor (n340, n308_mux, n311_mux);
xor (n340, n308, n311);
xnor (n340_xnor, n340, n340);
xor (n341, n340_mux, n315_mux);
xor (n341, n340, n315);
xnor (n341_xnor, n341, n341);
and (n342, n339_mux, n341_mux);
and (n342, n339, n341);
xnor (n342_xnor, n342, n342);
xor (n346, n343_mux, n345_mux);
xor (n346, n343, n345);
xnor (n346_xnor, n346, n346);
xor (n353, n346_mux, n352_mux);
xor (n353, n346, n352);
xnor (n353_xnor, n353, n353);
and (n354, n341_mux, n353_mux);
and (n354, n341, n353);
xnor (n354_xnor, n354, n354);
and (n355, n339_mux, n353_mux);
and (n355, n339, n353);
xnor (n355_xnor, n355, n355);
or (n356_1, n354_mux, n355_mux);
or (n356, n342_mux, n356_1);
or (n356_1, n354, n355);
or (n356, n342, n356_1);
xnor (n356_xnor, n356, n356);
and (n1310, n318_mux, n356_mux);
and (n1310, n318, n356);
xnor (n1310_xnor, n1310, n1310);
xor (n378, n361_mux, n377_mux);
xor (n378, n361, n377);
xnor (n378_xnor, n378, n378);
xor (n390, n378_mux, n389_mux);
xor (n390, n378, n389);
xnor (n390_xnor, n390, n390);
and (n1311, n356_mux, n390_mux);
and (n1311, n356, n390);
xnor (n1311_xnor, n1311, n1311);
and (n1312, n318_mux, n390_mux);
and (n1312, n318, n390);
xnor (n1312_xnor, n1312, n1312);
or (n1313_1, n1311_mux, n1312_mux);
or (n1313, n1310_mux, n1313_1);
or (n1313_1, n1311, n1312);
or (n1313, n1310, n1313_1);
xnor (n1313_xnor, n1313, n1313);
and (n1314, n1309_mux, n1313_mux);
and (n1314, n1309, n1313);
xnor (n1314_xnor, n1314, n1314);
xor (n1315, n1309_mux, n1313_mux);
xor (n1315, n1309, n1313);
xnor (n1315_xnor, n1315, n1315);
xor (n357, n318_mux, n356_mux);
xor (n357, n318, n356);
xnor (n357_xnor, n357, n357);
xor (n391, n357_mux, n390_mux);
xor (n391, n357, n390);
xnor (n391_xnor, n391, n391);
and (n392, n309_mux, n314_mux);
and (n392, n309, n314);
xnor (n392_xnor, n392, n392);
and (n393, n313_mux, n344_mux);
and (n393, n313, n344);
xnor (n393_xnor, n393, n393);
and (n394, n392_mux, n393_mux);
and (n394, n392, n393);
xnor (n394_xnor, n394, n394);
and (n395, n309_mux, n319_mux);
and (n395, n309, n319);
xnor (n395_xnor, n395, n395);
and (n396, n313_mux, n322_mux);
and (n396, n313, n322);
xnor (n396_xnor, n396, n396);
and (n397, n395_mux, n396_mux);
and (n397, n395, n396);
xnor (n397_xnor, n397, n397);
and (n398, n321_mux, n326_mux);
and (n398, n321, n326);
xnor (n398_xnor, n398, n398);
and (n399, n396_mux, n398_mux);
and (n399, n396, n398);
xnor (n399_xnor, n399, n399);
and (n400, n395_mux, n398_mux);
and (n400, n395, n398);
xnor (n400_xnor, n400, n400);
or (n401_1, n399_mux, n400_mux);
or (n401, n397_mux, n401_1);
or (n401_1, n399, n400);
or (n401, n397, n401_1);
xnor (n401_xnor, n401, n401);
and (n402, n309_mux, n344_mux);
and (n402, n309, n344);
xnor (n402_xnor, n402, n402);
and (n403, n401_mux, n402_mux);
and (n403, n401, n402);
xnor (n403_xnor, n403, n403);
xor (n404, n320_mux, n323_mux);
xor (n404, n320, n323);
xnor (n404_xnor, n404, n404);
xor (n405, n404_mux, n327_mux);
xor (n405, n404, n327);
xnor (n405_xnor, n405, n405);
and (n406, n402_mux, n405_mux);
and (n406, n402, n405);
xnor (n406_xnor, n406, n406);
and (n407, n401_mux, n405_mux);
and (n407, n401, n405);
xnor (n407_xnor, n407, n407);
or (n408_1, n406_mux, n407_mux);
or (n408, n403_mux, n408_1);
or (n408_1, n406, n407);
or (n408, n403, n408_1);
xnor (n408_xnor, n408, n408);
xor (n409, n392_mux, n393_mux);
xor (n409, n392, n393);
xnor (n409_xnor, n409, n409);
and (n410, n408_mux, n409_mux);
and (n410, n408, n409);
xnor (n410_xnor, n410, n410);
xor (n411, n330_mux, n331_mux);
xor (n411, n330, n331);
xnor (n411_xnor, n411, n411);
xor (n412, n411_mux, n336_mux);
xor (n412, n411, n336);
xnor (n412_xnor, n412, n412);
and (n413, n409_mux, n412_mux);
and (n413, n409, n412);
xnor (n413_xnor, n413, n413);
and (n414, n408_mux, n412_mux);
and (n414, n408, n412);
xnor (n414_xnor, n414, n414);
or (n415_1, n413_mux, n414_mux);
or (n415, n410_mux, n415_1);
or (n415_1, n413, n414);
or (n415, n410, n415_1);
xnor (n415_xnor, n415, n415);
and (n416, n394_mux, n415_mux);
and (n416, n394, n415);
xnor (n416_xnor, n416, n416);
xor (n417, n339_mux, n341_mux);
xor (n417, n339, n341);
xnor (n417_xnor, n417, n417);
xor (n418, n417_mux, n353_mux);
xor (n418, n417, n353);
xnor (n418_xnor, n418, n418);
and (n419, n415_mux, n418_mux);
and (n419, n415, n418);
xnor (n419_xnor, n419, n419);
and (n420, n394_mux, n418_mux);
and (n420, n394, n418);
xnor (n420_xnor, n420, n420);
or (n421_1, n419_mux, n420_mux);
or (n421, n416_mux, n421_1);
or (n421_1, n419, n420);
or (n421, n416, n421_1);
xnor (n421_xnor, n421, n421);
and (n1316, n391_mux, n421_mux);
and (n1316, n391, n421);
xnor (n1316_xnor, n1316, n1316);
xor (n422, n391_mux, n421_mux);
xor (n422, n391, n421);
xnor (n422_xnor, n422, n422);
xor (n423, n394_mux, n415_mux);
xor (n423, n394, n415);
xnor (n423_xnor, n423, n423);
xor (n424, n423_mux, n418_mux);
xor (n424, n423, n418);
xnor (n424_xnor, n424, n424);
and (n425, n306_mux, n319_mux);
and (n425, n306, n319);
xnor (n425_xnor, n425, n425);
and (n426, n309_mux, n322_mux);
and (n426, n309, n322);
xnor (n426_xnor, n426, n426);
and (n427, n425_mux, n426_mux);
and (n427, n425, n426);
xnor (n427_xnor, n427, n427);
and (n428, n313_mux, n326_mux);
and (n428, n313, n326);
xnor (n428_xnor, n428, n428);
and (n429, n426_mux, n428_mux);
and (n429, n426, n428);
xnor (n429_xnor, n429, n429);
and (n430, n425_mux, n428_mux);
and (n430, n425, n428);
xnor (n430_xnor, n430, n430);
or (n431_1, n429_mux, n430_mux);
or (n431, n427_mux, n431_1);
or (n431_1, n429, n430);
or (n431, n427, n431_1);
xnor (n431_xnor, n431, n431);
and (n432, n306_mux, n344_mux);
and (n432, n306, n344);
xnor (n432_xnor, n432, n432);
and (n433, n431_mux, n432_mux);
and (n433, n431, n432);
xnor (n433_xnor, n433, n433);
xor (n434, n395_mux, n396_mux);
xor (n434, n395, n396);
xnor (n434_xnor, n434, n434);
xor (n435, n434_mux, n398_mux);
xor (n435, n434, n398);
xnor (n435_xnor, n435, n435);
and (n436, n432_mux, n435_mux);
and (n436, n432, n435);
xnor (n436_xnor, n436, n436);
and (n437, n431_mux, n435_mux);
and (n437, n431, n435);
xnor (n437_xnor, n437, n437);
or (n438_1, n436_mux, n437_mux);
or (n438, n433_mux, n438_1);
or (n438_1, n436, n437);
or (n438, n433, n438_1);
xnor (n438_xnor, n438, n438);
and (n439, n306_mux, n314_mux);
and (n439, n306, n314);
xnor (n439_xnor, n439, n439);
and (n440, n438_mux, n439_mux);
and (n440, n438, n439);
xnor (n440_xnor, n440, n440);
xor (n441, n401_mux, n402_mux);
xor (n441, n401, n402);
xnor (n441_xnor, n441, n441);
xor (n442, n441_mux, n405_mux);
xor (n442, n441, n405);
xnor (n442_xnor, n442, n442);
and (n443, n439_mux, n442_mux);
and (n443, n439, n442);
xnor (n443_xnor, n443, n443);
and (n444, n438_mux, n442_mux);
and (n444, n438, n442);
xnor (n444_xnor, n444, n444);
or (n445_1, n443_mux, n444_mux);
or (n445, n440_mux, n445_1);
or (n445_1, n443, n444);
or (n445, n440, n445_1);
xnor (n445_xnor, n445, n445);
xor (n446, n408_mux, n409_mux);
xor (n446, n408, n409);
xnor (n446_xnor, n446, n446);
xor (n447, n446_mux, n412_mux);
xor (n447, n446, n412);
xnor (n447_xnor, n447, n447);
and (n448, n445_mux, n447_mux);
and (n448, n445, n447);
xnor (n448_xnor, n448, n448);
and (n449, n424_mux, n448_mux);
and (n449, n424, n448);
xnor (n449_xnor, n449, n449);
xor (n450, n424_mux, n448_mux);
xor (n450, n424, n448);
xnor (n450_xnor, n450, n450);
and (n451, n306_mux, n310_mux);
and (n451, n306, n310);
xnor (n451_xnor, n451, n451);
xor (n452, n445_mux, n447_mux);
xor (n452, n445, n447);
xnor (n452_xnor, n452, n452);
and (n453, n451_mux, n452_mux);
and (n453, n451, n452);
xnor (n453_xnor, n453, n453);
xor (n454, n451_mux, n452_mux);
xor (n454, n451, n452);
xnor (n454_xnor, n454, n454);
xor (n455, n438_mux, n439_mux);
xor (n455, n438, n439);
xnor (n455_xnor, n455, n455);
xor (n456, n455_mux, n442_mux);
xor (n456, n455, n442);
xnor (n456_xnor, n456, n456);
xor (n457, n431_mux, n432_mux);
xor (n457, n431, n432);
xnor (n457_xnor, n457, n457);
xor (n458, n457_mux, n435_mux);
xor (n458, n457, n435);
xnor (n458_xnor, n458, n458);
xor (n459, n425_mux, n426_mux);
xor (n459, n425, n426);
xnor (n459_xnor, n459, n459);
xor (n460, n459_mux, n428_mux);
xor (n460, n459, n428);
xnor (n460_xnor, n460, n460);
and (n461, n306_mux, n322_mux);
and (n461, n306, n322);
xnor (n461_xnor, n461, n461);
and (n462, n309_mux, n326_mux);
and (n462, n309, n326);
xnor (n462_xnor, n462, n462);
and (n463, n461_mux, n462_mux);
and (n463, n461, n462);
xnor (n463_xnor, n463, n463);
and (n464, n460_mux, n463_mux);
and (n464, n460, n463);
xnor (n464_xnor, n464, n464);
and (n465, n458_mux, n464_mux);
and (n465, n458, n464);
xnor (n465_xnor, n465, n465);
and (n466, n456_mux, n465_mux);
and (n466, n456, n465);
xnor (n466_xnor, n466, n466);
and (n467, n454_mux, n466_mux);
and (n467, n454, n466);
xnor (n467_xnor, n467, n467);
or (n468, n453_mux, n467_mux);
or (n468, n453, n467);
xnor (n468_xnor, n468, n468);
and (n469, n450_mux, n468_mux);
and (n469, n450, n468);
xnor (n469_xnor, n469, n469);
or (n470, n449_mux, n469_mux);
or (n470, n449, n469);
xnor (n470_xnor, n470, n470);
and (n1317, n422_mux, n470_mux);
and (n1317, n422, n470);
xnor (n1317_xnor, n1317, n1317);
or (n1318, n1316_mux, n1317_mux);
or (n1318, n1316, n1317);
xnor (n1318_xnor, n1318, n1318);
and (n1319, n1315_mux, n1318_mux);
and (n1319, n1315, n1318);
xnor (n1319_xnor, n1319, n1319);
or (n1320, n1314_mux, n1319_mux);
or (n1320, n1314, n1319);
xnor (n1320_xnor, n1320, n1320);
and (n1321, n1307_mux, n1320_mux);
and (n1321, n1307, n1320);
xnor (n1321_xnor, n1321, n1321);
or (n1322, n1306_mux, n1321_mux);
or (n1322, n1306, n1321);
xnor (n1322_xnor, n1322, n1322);
and (n1323, n1292_mux, n1322_mux);
and (n1323, n1292, n1322);
xnor (n1323_xnor, n1323, n1323);
or (n1324, n1291_mux, n1323_mux);
or (n1324, n1291, n1323);
xnor (n1324_xnor, n1324, n1324);
and (n1325, n1256_mux, n1324_mux);
and (n1325, n1256, n1324);
xnor (n1325_xnor, n1325, n1325);
or (n1326, n1255_mux, n1325_mux);
or (n1326, n1255, n1325);
xnor (n1326_xnor, n1326, n1326);
and (n1327, n1216_mux, n1326_mux);
and (n1327, n1216, n1326);
xnor (n1327_xnor, n1327, n1327);
or (n1328, n1215_mux, n1327_mux);
or (n1328, n1215, n1327);
xnor (n1328_xnor, n1328, n1328);
and (n1329, n1179_mux, n1328_mux);
and (n1329, n1179, n1328);
xnor (n1329_xnor, n1329, n1329);
or (n1330, n1178_mux, n1329_mux);
or (n1330, n1178, n1329);
xnor (n1330_xnor, n1330, n1330);
and (n1331, n1136_mux, n1330_mux);
and (n1331, n1136, n1330);
xnor (n1331_xnor, n1331, n1331);
or (n1332, n1135_mux, n1331_mux);
or (n1332, n1135, n1331);
xnor (n1332_xnor, n1332, n1332);
buf(n1333, n1332_mux);
buf(n1333, n1332);
xnor (n1333_xnor, n1333, n1333);
buf(n1463, n1333_mux);
buf(n1463, n1333);
xnor (n1463_xnor, n1463, n1463);
xor (n1334, n1136_mux, n1330_mux);
xor (n1334, n1136, n1330);
xnor (n1334_xnor, n1334, n1334);
buf(n1335, n1334_mux);
buf(n1335, n1334);
xnor (n1335_xnor, n1335, n1335);
buf(n1464, n1335_mux);
buf(n1464, n1335);
xnor (n1464_xnor, n1464, n1464);
xor (n1336, n1179_mux, n1328_mux);
xor (n1336, n1179, n1328);
xnor (n1336_xnor, n1336, n1336);
buf(n1337, n1336_mux);
buf(n1337, n1336);
xnor (n1337_xnor, n1337, n1337);
buf(n1465, n1337_mux);
buf(n1465, n1337);
xnor (n1465_xnor, n1465, n1465);
xor (n1338, n1216_mux, n1326_mux);
xor (n1338, n1216, n1326);
xnor (n1338_xnor, n1338, n1338);
buf(n1339, n1338_mux);
buf(n1339, n1338);
xnor (n1339_xnor, n1339, n1339);
buf(n1466, n1339_mux);
buf(n1466, n1339);
xnor (n1466_xnor, n1466, n1466);
xor (n1340, n1256_mux, n1324_mux);
xor (n1340, n1256, n1324);
xnor (n1340_xnor, n1340, n1340);
buf(n1341, n1340_mux);
buf(n1341, n1340);
xnor (n1341_xnor, n1341, n1341);
buf(n1467, n1341_mux);
buf(n1467, n1341);
xnor (n1467_xnor, n1467, n1467);
xor (n1342, n1292_mux, n1322_mux);
xor (n1342, n1292, n1322);
xnor (n1342_xnor, n1342, n1342);
buf(n1343, n1342_mux);
buf(n1343, n1342);
xnor (n1343_xnor, n1343, n1343);
buf(n1468, n1343_mux);
buf(n1468, n1343);
xnor (n1468_xnor, n1468, n1468);
xor (n1344, n1307_mux, n1320_mux);
xor (n1344, n1307, n1320);
xnor (n1344_xnor, n1344, n1344);
buf(n1345, n1344_mux);
buf(n1345, n1344);
xnor (n1345_xnor, n1345, n1345);
buf(n1469, n1345_mux);
buf(n1469, n1345);
xnor (n1469_xnor, n1469, n1469);
xor (n638, n450_mux, n468_mux);
xor (n638, n450, n468);
xnor (n638_xnor, n638, n638);
buf(n639, n638_mux);
buf(n639, n638);
xnor (n639_xnor, n639, n639);
buf(n640, n639_mux);
buf(n640, n639);
xnor (n640_xnor, n640, n640);
xnor (g14_xnor, g14, g14);
buf(n33, g14_mux);
buf(n33, g14);
xnor (n33_xnor, n33, n33);
buf(n474, n33_mux);
buf(n474, n33);
xnor (n474_xnor, n474, n474);
xnor (g27_xnor, g27, g27);
buf(n46, g27_mux);
buf(n46, g27);
xnor (n46_xnor, n46, n46);
buf(n479, n46_mux);
buf(n479, n46);
xnor (n479_xnor, n479, n479);
and (n557, n474_mux, n479_mux);
and (n557, n474, n479);
xnor (n557_xnor, n557, n557);
xnor (g13_xnor, g13, g13);
buf(n32, g13_mux);
buf(n32, g13);
xnor (n32_xnor, n32, n32);
buf(n478, n32_mux);
buf(n478, n32);
xnor (n478_xnor, n478, n478);
xnor (g28_xnor, g28, g28);
buf(n47, g28_mux);
buf(n47, g28);
xnor (n47_xnor, n47, n47);
buf(n509, n47_mux);
buf(n509, n47);
xnor (n509_xnor, n509, n509);
and (n558, n478_mux, n509_mux);
and (n558, n478, n509);
xnor (n558_xnor, n558, n558);
and (n559, n557_mux, n558_mux);
and (n559, n557, n558);
xnor (n559_xnor, n559, n559);
xnor (g29_xnor, g29, g29);
buf(n48, g29_mux);
buf(n48, g29);
xnor (n48_xnor, n48, n48);
buf(n484, n48_mux);
buf(n484, n48);
xnor (n484_xnor, n484, n484);
and (n560, n474_mux, n484_mux);
and (n560, n474, n484);
xnor (n560_xnor, n560, n560);
xnor (g30_xnor, g30, g30);
buf(n49, g30_mux);
buf(n49, g30);
xnor (n49_xnor, n49, n49);
buf(n487, n49_mux);
buf(n487, n49);
xnor (n487_xnor, n487, n487);
and (n561, n478_mux, n487_mux);
and (n561, n478, n487);
xnor (n561_xnor, n561, n561);
and (n562, n560_mux, n561_mux);
and (n562, n560, n561);
xnor (n562_xnor, n562, n562);
xnor (g12_xnor, g12, g12);
buf(n31, g12_mux);
buf(n31, g12);
xnor (n31_xnor, n31, n31);
buf(n486, n31_mux);
buf(n486, n31);
xnor (n486_xnor, n486, n486);
xnor (g31_xnor, g31, g31);
buf(n50, g31_mux);
buf(n50, g31);
xnor (n50_xnor, n50, n50);
buf(n491, n50_mux);
buf(n491, n50);
xnor (n491_xnor, n491, n491);
and (n563, n486_mux, n491_mux);
and (n563, n486, n491);
xnor (n563_xnor, n563, n563);
and (n564, n561_mux, n563_mux);
and (n564, n561, n563);
xnor (n564_xnor, n564, n564);
and (n565, n560_mux, n563_mux);
and (n565, n560, n563);
xnor (n565_xnor, n565, n565);
or (n566_1, n564_mux, n565_mux);
or (n566, n562_mux, n566_1);
or (n566_1, n564, n565);
or (n566, n562, n566_1);
xnor (n566_xnor, n566, n566);
and (n567, n474_mux, n509_mux);
and (n567, n474, n509);
xnor (n567_xnor, n567, n567);
and (n568, n566_mux, n567_mux);
and (n568, n566, n567);
xnor (n568_xnor, n568, n568);
and (n485, n478_mux, n484_mux);
and (n485, n478, n484);
xnor (n485_xnor, n485, n485);
and (n488, n486_mux, n487_mux);
and (n488, n486, n487);
xnor (n488_xnor, n488, n488);
xor (n569, n485_mux, n488_mux);
xor (n569, n485, n488);
xnor (n569_xnor, n569, n569);
xnor (g11_xnor, g11, g11);
buf(n30, g11_mux);
buf(n30, g11);
xnor (n30_xnor, n30, n30);
buf(n490, n30_mux);
buf(n490, n30);
xnor (n490_xnor, n490, n490);
and (n492, n490_mux, n491_mux);
and (n492, n490, n491);
xnor (n492_xnor, n492, n492);
xor (n570, n569_mux, n492_mux);
xor (n570, n569, n492);
xnor (n570_xnor, n570, n570);
and (n571, n567_mux, n570_mux);
and (n571, n567, n570);
xnor (n571_xnor, n571, n571);
and (n572, n566_mux, n570_mux);
and (n572, n566, n570);
xnor (n572_xnor, n572, n572);
or (n573_1, n571_mux, n572_mux);
or (n573, n568_mux, n573_1);
or (n573_1, n571, n572);
or (n573, n568, n573_1);
xnor (n573_xnor, n573, n573);
xor (n574, n557_mux, n558_mux);
xor (n574, n557, n558);
xnor (n574_xnor, n574, n574);
and (n575, n573_mux, n574_mux);
and (n575, n573, n574);
xnor (n575_xnor, n575, n575);
and (n489, n485_mux, n488_mux);
and (n489, n485, n488);
xnor (n489_xnor, n489, n489);
and (n493, n488_mux, n492_mux);
and (n493, n488, n492);
xnor (n493_xnor, n493, n493);
and (n494, n485_mux, n492_mux);
and (n494, n485, n492);
xnor (n494_xnor, n494, n494);
or (n495_1, n493_mux, n494_mux);
or (n495, n489_mux, n495_1);
or (n495_1, n493, n494);
or (n495, n489, n495_1);
xnor (n495_xnor, n495, n495);
and (n496, n486_mux, n484_mux);
and (n496, n486, n484);
xnor (n496_xnor, n496, n496);
xor (n576, n495_mux, n496_mux);
xor (n576, n495, n496);
xnor (n576_xnor, n576, n576);
and (n498, n490_mux, n487_mux);
and (n498, n490, n487);
xnor (n498_xnor, n498, n498);
xnor (g10_xnor, g10, g10);
buf(n29, g10_mux);
buf(n29, g10);
xnor (n29_xnor, n29, n29);
buf(n499, n29_mux);
buf(n499, n29);
xnor (n499_xnor, n499, n499);
and (n500, n499_mux, n491_mux);
and (n500, n499, n491);
xnor (n500_xnor, n500, n500);
xor (n501, n498_mux, n500_mux);
xor (n501, n498, n500);
xnor (n501_xnor, n501, n501);
xor (n577, n576_mux, n501_mux);
xor (n577, n576, n501);
xnor (n577_xnor, n577, n577);
and (n578, n574_mux, n577_mux);
and (n578, n574, n577);
xnor (n578_xnor, n578, n578);
and (n579, n573_mux, n577_mux);
and (n579, n573, n577);
xnor (n579_xnor, n579, n579);
or (n580_1, n578_mux, n579_mux);
or (n580, n575_mux, n580_1);
or (n580_1, n578, n579);
or (n580, n575, n580_1);
xnor (n580_xnor, n580, n580);
xor (n588, n559_mux, n580_mux);
xor (n588, n559, n580);
xnor (n588_xnor, n588, n588);
and (n497, n495_mux, n496_mux);
and (n497, n495, n496);
xnor (n497_xnor, n497, n497);
and (n502, n496_mux, n501_mux);
and (n502, n496, n501);
xnor (n502_xnor, n502, n502);
and (n503, n495_mux, n501_mux);
and (n503, n495, n501);
xnor (n503_xnor, n503, n503);
or (n504_1, n502_mux, n503_mux);
or (n504, n497_mux, n504_1);
or (n504_1, n502, n503);
or (n504, n497, n504_1);
xnor (n504_xnor, n504, n504);
xnor (g15_xnor, g15, g15);
buf(n34, g15_mux);
buf(n34, g15);
xnor (n34_xnor, n34, n34);
buf(n471, n34_mux);
buf(n471, n34);
xnor (n471_xnor, n471, n471);
xnor (g25_xnor, g25, g25);
buf(n44, g25_mux);
buf(n44, g25);
xnor (n44_xnor, n44, n44);
buf(n472, n44_mux);
buf(n472, n44);
xnor (n472_xnor, n472, n472);
and (n473, n471_mux, n472_mux);
and (n473, n471, n472);
xnor (n473_xnor, n473, n473);
xnor (g26_xnor, g26, g26);
buf(n45, g26_mux);
buf(n45, g26);
xnor (n45_xnor, n45, n45);
buf(n475, n45_mux);
buf(n475, n45);
xnor (n475_xnor, n475, n475);
and (n476, n474_mux, n475_mux);
and (n476, n474, n475);
xnor (n476_xnor, n476, n476);
xor (n505, n473_mux, n476_mux);
xor (n505, n473, n476);
xnor (n505_xnor, n505, n505);
and (n480, n478_mux, n479_mux);
and (n480, n478, n479);
xnor (n480_xnor, n480, n480);
xor (n506, n505_mux, n480_mux);
xor (n506, n505, n480);
xnor (n506_xnor, n506, n506);
xor (n582, n504_mux, n506_mux);
xor (n582, n504, n506);
xnor (n582_xnor, n582, n582);
and (n508, n498_mux, n500_mux);
and (n508, n498, n500);
xnor (n508_xnor, n508, n508);
and (n510, n486_mux, n509_mux);
and (n510, n486, n509);
xnor (n510_xnor, n510, n510);
xor (n511, n508_mux, n510_mux);
xor (n511, n508, n510);
xnor (n511_xnor, n511, n511);
and (n512, n490_mux, n484_mux);
and (n512, n490, n484);
xnor (n512_xnor, n512, n512);
and (n513, n499_mux, n487_mux);
and (n513, n499, n487);
xnor (n513_xnor, n513, n513);
xor (n514, n512_mux, n513_mux);
xor (n514, n512, n513);
xnor (n514_xnor, n514, n514);
xnor (g9_xnor, g9, g9);
buf(n28, g9_mux);
buf(n28, g9);
xnor (n28_xnor, n28, n28);
buf(n515, n28_mux);
buf(n515, n28);
xnor (n515_xnor, n515, n515);
and (n516, n515_mux, n491_mux);
and (n516, n515, n491);
xnor (n516_xnor, n516, n516);
xor (n517, n514_mux, n516_mux);
xor (n517, n514, n516);
xnor (n517_xnor, n517, n517);
xor (n518, n511_mux, n517_mux);
xor (n518, n511, n517);
xnor (n518_xnor, n518, n518);
xor (n583, n582_mux, n518_mux);
xor (n583, n582, n518);
xnor (n583_xnor, n583, n583);
xor (n589, n588_mux, n583_mux);
xor (n589, n588, n583);
xnor (n589_xnor, n589, n589);
and (n590, n471_mux, n484_mux);
and (n590, n471, n484);
xnor (n590_xnor, n590, n590);
and (n591, n474_mux, n487_mux);
and (n591, n474, n487);
xnor (n591_xnor, n591, n591);
and (n592, n590_mux, n591_mux);
and (n592, n590, n591);
xnor (n592_xnor, n592, n592);
and (n593, n478_mux, n491_mux);
and (n593, n478, n491);
xnor (n593_xnor, n593, n593);
and (n594, n591_mux, n593_mux);
and (n594, n591, n593);
xnor (n594_xnor, n594, n594);
and (n595, n590_mux, n593_mux);
and (n595, n590, n593);
xnor (n595_xnor, n595, n595);
or (n596_1, n594_mux, n595_mux);
or (n596, n592_mux, n596_1);
or (n596_1, n594, n595);
or (n596, n592, n596_1);
xnor (n596_xnor, n596, n596);
and (n597, n471_mux, n509_mux);
and (n597, n471, n509);
xnor (n597_xnor, n597, n597);
and (n598, n596_mux, n597_mux);
and (n598, n596, n597);
xnor (n598_xnor, n598, n598);
xor (n599, n560_mux, n561_mux);
xor (n599, n560, n561);
xnor (n599_xnor, n599, n599);
xor (n600, n599_mux, n563_mux);
xor (n600, n599, n563);
xnor (n600_xnor, n600, n600);
and (n601, n597_mux, n600_mux);
and (n601, n597, n600);
xnor (n601_xnor, n601, n601);
and (n602, n596_mux, n600_mux);
and (n602, n596, n600);
xnor (n602_xnor, n602, n602);
or (n603_1, n601_mux, n602_mux);
or (n603, n598_mux, n603_1);
or (n603_1, n601, n602);
or (n603, n598, n603_1);
xnor (n603_xnor, n603, n603);
and (n604, n471_mux, n479_mux);
and (n604, n471, n479);
xnor (n604_xnor, n604, n604);
and (n605, n603_mux, n604_mux);
and (n605, n603, n604);
xnor (n605_xnor, n605, n605);
xor (n606, n566_mux, n567_mux);
xor (n606, n566, n567);
xnor (n606_xnor, n606, n606);
xor (n607, n606_mux, n570_mux);
xor (n607, n606, n570);
xnor (n607_xnor, n607, n607);
and (n608, n604_mux, n607_mux);
and (n608, n604, n607);
xnor (n608_xnor, n608, n608);
and (n609, n603_mux, n607_mux);
and (n609, n603, n607);
xnor (n609_xnor, n609, n609);
or (n610_1, n608_mux, n609_mux);
or (n610, n605_mux, n610_1);
or (n610_1, n608, n609);
or (n610, n605, n610_1);
xnor (n610_xnor, n610, n610);
xor (n611, n573_mux, n574_mux);
xor (n611, n573, n574);
xnor (n611_xnor, n611, n611);
xor (n612, n611_mux, n577_mux);
xor (n612, n611, n577);
xnor (n612_xnor, n612, n612);
and (n613, n610_mux, n612_mux);
and (n613, n610, n612);
xnor (n613_xnor, n613, n613);
xor (n615, n589_mux, n613_mux);
xor (n615, n589, n613);
xnor (n615_xnor, n615, n615);
and (n616, n471_mux, n475_mux);
and (n616, n471, n475);
xnor (n616_xnor, n616, n616);
xor (n617, n610_mux, n612_mux);
xor (n617, n610, n612);
xnor (n617_xnor, n617, n617);
and (n618, n616_mux, n617_mux);
and (n618, n616, n617);
xnor (n618_xnor, n618, n618);
xor (n619, n616_mux, n617_mux);
xor (n619, n616, n617);
xnor (n619_xnor, n619, n619);
xor (n620, n603_mux, n604_mux);
xor (n620, n603, n604);
xnor (n620_xnor, n620, n620);
xor (n621, n620_mux, n607_mux);
xor (n621, n620, n607);
xnor (n621_xnor, n621, n621);
xor (n622, n596_mux, n597_mux);
xor (n622, n596, n597);
xnor (n622_xnor, n622, n622);
xor (n623, n622_mux, n600_mux);
xor (n623, n622, n600);
xnor (n623_xnor, n623, n623);
xor (n624, n590_mux, n591_mux);
xor (n624, n590, n591);
xnor (n624_xnor, n624, n624);
xor (n625, n624_mux, n593_mux);
xor (n625, n624, n593);
xnor (n625_xnor, n625, n625);
and (n626, n471_mux, n487_mux);
and (n626, n471, n487);
xnor (n626_xnor, n626, n626);
and (n627, n474_mux, n491_mux);
and (n627, n474, n491);
xnor (n627_xnor, n627, n627);
and (n628, n626_mux, n627_mux);
and (n628, n626, n627);
xnor (n628_xnor, n628, n628);
and (n629, n625_mux, n628_mux);
and (n629, n625, n628);
xnor (n629_xnor, n629, n629);
and (n630, n623_mux, n629_mux);
and (n630, n623, n629);
xnor (n630_xnor, n630, n630);
and (n631, n621_mux, n630_mux);
and (n631, n621, n630);
xnor (n631_xnor, n631, n631);
and (n632, n619_mux, n631_mux);
and (n632, n619, n631);
xnor (n632_xnor, n632, n632);
or (n633, n618_mux, n632_mux);
or (n633, n618, n632);
xnor (n633_xnor, n633, n633);
xor (n641, n615_mux, n633_mux);
xor (n641, n615, n633);
xnor (n641_xnor, n641, n641);
buf(n642, n641_mux);
buf(n642, n641);
xnor (n642_xnor, n642, n642);
buf(n643, n642_mux);
buf(n643, n642);
xnor (n643_xnor, n643, n643);
and (n644, n640_mux, n643_mux);
and (n644, n640, n643);
xnor (n644_xnor, n644, n644);
xor (n645, n454_mux, n466_mux);
xor (n645, n454, n466);
xnor (n645_xnor, n645, n645);
buf(n646, n645_mux);
buf(n646, n645);
xnor (n646_xnor, n646, n646);
buf(n647, n646_mux);
buf(n647, n646);
xnor (n647_xnor, n647, n647);
xor (n648, n619_mux, n631_mux);
xor (n648, n619, n631);
xnor (n648_xnor, n648, n648);
buf(n649, n648_mux);
buf(n649, n648);
xnor (n649_xnor, n649, n649);
buf(n650, n649_mux);
buf(n650, n649);
xnor (n650_xnor, n650, n650);
and (n651, n647_mux, n650_mux);
and (n651, n647, n650);
xnor (n651_xnor, n651, n651);
xor (n652, n456_mux, n465_mux);
xor (n652, n456, n465);
xnor (n652_xnor, n652, n652);
buf(n653, n652_mux);
buf(n653, n652);
xnor (n653_xnor, n653, n653);
buf(n654, n653_mux);
buf(n654, n653);
xnor (n654_xnor, n654, n654);
xor (n655, n621_mux, n630_mux);
xor (n655, n621, n630);
xnor (n655_xnor, n655, n655);
buf(n656, n655_mux);
buf(n656, n655);
xnor (n656_xnor, n656, n656);
buf(n657, n656_mux);
buf(n657, n656);
xnor (n657_xnor, n657, n657);
and (n658, n654_mux, n657_mux);
and (n658, n654, n657);
xnor (n658_xnor, n658, n658);
xor (n659, n458_mux, n464_mux);
xor (n659, n458, n464);
xnor (n659_xnor, n659, n659);
buf(n660, n659_mux);
buf(n660, n659);
xnor (n660_xnor, n660, n660);
buf(n661, n660_mux);
buf(n661, n660);
xnor (n661_xnor, n661, n661);
xor (n662, n623_mux, n629_mux);
xor (n662, n623, n629);
xnor (n662_xnor, n662, n662);
buf(n663, n662_mux);
buf(n663, n662);
xnor (n663_xnor, n663, n663);
buf(n664, n663_mux);
buf(n664, n663);
xnor (n664_xnor, n664, n664);
and (n665, n661_mux, n664_mux);
and (n665, n661, n664);
xnor (n665_xnor, n665, n665);
xor (n666, n460_mux, n463_mux);
xor (n666, n460, n463);
xnor (n666_xnor, n666, n666);
buf(n667, n666_mux);
buf(n667, n666);
xnor (n667_xnor, n667, n667);
buf(n668, n667_mux);
buf(n668, n667);
xnor (n668_xnor, n668, n668);
xor (n669, n625_mux, n628_mux);
xor (n669, n625, n628);
xnor (n669_xnor, n669, n669);
buf(n670, n669_mux);
buf(n670, n669);
xnor (n670_xnor, n670, n670);
buf(n671, n670_mux);
buf(n671, n670);
xnor (n671_xnor, n671, n671);
and (n672, n668_mux, n671_mux);
and (n672, n668, n671);
xnor (n672_xnor, n672, n672);
xor (n673, n461_mux, n462_mux);
xor (n673, n461, n462);
xnor (n673_xnor, n673, n673);
buf(n674, n673_mux);
buf(n674, n673);
xnor (n674_xnor, n674, n674);
buf(n675, n674_mux);
buf(n675, n674);
xnor (n675_xnor, n675, n675);
xor (n676, n626_mux, n627_mux);
xor (n676, n626, n627);
xnor (n676_xnor, n676, n676);
buf(n677, n676_mux);
buf(n677, n676);
xnor (n677_xnor, n677, n677);
buf(n678, n677_mux);
buf(n678, n677);
xnor (n678_xnor, n678, n678);
and (n679, n675_mux, n678_mux);
and (n679, n675, n678);
xnor (n679_xnor, n679, n679);
and (n680, n306_mux, n326_mux);
and (n680, n306, n326);
xnor (n680_xnor, n680, n680);
buf(n681, n680_mux);
buf(n681, n680);
xnor (n681_xnor, n681, n681);
buf(n682, n681_mux);
buf(n682, n681);
xnor (n682_xnor, n682, n682);
and (n683, n471_mux, n491_mux);
and (n683, n471, n491);
xnor (n683_xnor, n683, n683);
buf(n684, n683_mux);
buf(n684, n683);
xnor (n684_xnor, n684, n684);
buf(n685, n684_mux);
buf(n685, n684);
xnor (n685_xnor, n685, n685);
and (n686, n682_mux, n685_mux);
and (n686, n682, n685);
xnor (n686_xnor, n686, n686);
and (n687, n678_mux, n686_mux);
and (n687, n678, n686);
xnor (n687_xnor, n687, n687);
and (n688, n675_mux, n686_mux);
and (n688, n675, n686);
xnor (n688_xnor, n688, n688);
or (n689_1, n687_mux, n688_mux);
or (n689, n679_mux, n689_1);
or (n689_1, n687, n688);
or (n689, n679, n689_1);
xnor (n689_xnor, n689, n689);
and (n690, n671_mux, n689_mux);
and (n690, n671, n689);
xnor (n690_xnor, n690, n690);
and (n691, n668_mux, n689_mux);
and (n691, n668, n689);
xnor (n691_xnor, n691, n691);
or (n692_1, n690_mux, n691_mux);
or (n692, n672_mux, n692_1);
or (n692_1, n690, n691);
or (n692, n672, n692_1);
xnor (n692_xnor, n692, n692);
and (n693, n664_mux, n692_mux);
and (n693, n664, n692);
xnor (n693_xnor, n693, n693);
and (n694, n661_mux, n692_mux);
and (n694, n661, n692);
xnor (n694_xnor, n694, n694);
or (n695_1, n693_mux, n694_mux);
or (n695, n665_mux, n695_1);
or (n695_1, n693, n694);
or (n695, n665, n695_1);
xnor (n695_xnor, n695, n695);
and (n696, n657_mux, n695_mux);
and (n696, n657, n695);
xnor (n696_xnor, n696, n696);
and (n697, n654_mux, n695_mux);
and (n697, n654, n695);
xnor (n697_xnor, n697, n697);
or (n698_1, n696_mux, n697_mux);
or (n698, n658_mux, n698_1);
or (n698_1, n696, n697);
or (n698, n658, n698_1);
xnor (n698_xnor, n698, n698);
and (n699, n650_mux, n698_mux);
and (n699, n650, n698);
xnor (n699_xnor, n699, n699);
and (n700, n647_mux, n698_mux);
and (n700, n647, n698);
xnor (n700_xnor, n700, n700);
or (n701_1, n699_mux, n700_mux);
or (n701, n651_mux, n701_1);
or (n701_1, n699, n700);
or (n701, n651, n701_1);
xnor (n701_xnor, n701, n701);
and (n702, n643_mux, n701_mux);
and (n702, n643, n701);
xnor (n702_xnor, n702, n702);
and (n703, n640_mux, n701_mux);
and (n703, n640, n701);
xnor (n703_xnor, n703, n703);
or (n704_1, n702_mux, n703_mux);
or (n704, n644_mux, n704_1);
or (n704_1, n702, n703);
or (n704, n644, n704_1);
xnor (n704_xnor, n704, n704);
xor (n705, t_0, n704_mux);
xor (n705, t_0, n704);
xnor (n705_xnor, n705, n705);
buf(n706, n705_mux);
buf(n706, n705);
xnor (n706_xnor, n706, n706);
not(n25, n706_mux);
not(n25, n706);
xnor (n25_xnor, n25, n25);
buf(n816, n35_mux);
buf(n816, n35);
xnor (n816_xnor, n816, n816);
xnor (g24_xnor, g24, g24);
buf(n43, g24_mux);
buf(n43, g24);
xnor (n43_xnor, n43, n43);
buf(n817, n43_mux);
buf(n817, n43);
xnor (n817_xnor, n817, n817);
and (n835, n816_mux, n817_mux);
and (n835, n816, n817);
xnor (n835_xnor, n835, n835);
buf(n797, n36_mux);
buf(n797, n36);
xnor (n797_xnor, n797, n797);
buf(n798, n44_mux);
buf(n798, n44);
xnor (n798_xnor, n798, n798);
and (n819, n797_mux, n798_mux);
and (n819, n797, n798);
xnor (n819_xnor, n819, n819);
buf(n778, n37_mux);
buf(n778, n37);
xnor (n778_xnor, n778, n778);
buf(n779, n45_mux);
buf(n779, n45);
xnor (n779_xnor, n779, n779);
and (n800, n778_mux, n779_mux);
and (n800, n778, n779);
xnor (n800_xnor, n800, n800);
buf(n759, n38_mux);
buf(n759, n38);
xnor (n759_xnor, n759, n759);
buf(n760, n46_mux);
buf(n760, n46);
xnor (n760_xnor, n760, n760);
and (n781, n759_mux, n760_mux);
and (n781, n759, n760);
xnor (n781_xnor, n781, n781);
buf(n740, n39_mux);
buf(n740, n39);
xnor (n740_xnor, n740, n740);
buf(n741, n47_mux);
buf(n741, n47);
xnor (n741_xnor, n741, n741);
and (n762, n740_mux, n741_mux);
and (n762, n740, n741);
xnor (n762_xnor, n762, n762);
buf(n721, n40_mux);
buf(n721, n40);
xnor (n721_xnor, n721, n721);
buf(n722, n48_mux);
buf(n722, n48);
xnor (n722_xnor, n722, n722);
and (n743, n721_mux, n722_mux);
and (n743, n721, n722);
xnor (n743_xnor, n743, n743);
buf(n708, n41_mux);
buf(n708, n41);
xnor (n708_xnor, n708, n708);
buf(n709, n49_mux);
buf(n709, n49);
xnor (n709_xnor, n709, n709);
and (n724, n708_mux, n709_mux);
and (n724, n708, n709);
xnor (n724_xnor, n724, n724);
buf(n298, n42_mux);
buf(n298, n42);
xnor (n298_xnor, n298, n298);
buf(n299, n50_mux);
buf(n299, n50);
xnor (n299_xnor, n299, n299);
and (n711, n298_mux, n299_mux);
and (n711, n298, n299);
xnor (n711_xnor, n711, n711);
and (n725, n709_mux, n711_mux);
and (n725, n709, n711);
xnor (n725_xnor, n725, n725);
and (n726, n708_mux, n711_mux);
and (n726, n708, n711);
xnor (n726_xnor, n726, n726);
or (n727_1, n725_mux, n726_mux);
or (n727, n724_mux, n727_1);
or (n727_1, n725, n726);
or (n727, n724, n727_1);
xnor (n727_xnor, n727, n727);
and (n744, n722_mux, n727_mux);
and (n744, n722, n727);
xnor (n744_xnor, n744, n744);
and (n745, n721_mux, n727_mux);
and (n745, n721, n727);
xnor (n745_xnor, n745, n745);
or (n746_1, n744_mux, n745_mux);
or (n746, n743_mux, n746_1);
or (n746_1, n744, n745);
or (n746, n743, n746_1);
xnor (n746_xnor, n746, n746);
and (n763, n741_mux, n746_mux);
and (n763, n741, n746);
xnor (n763_xnor, n763, n763);
and (n764, n740_mux, n746_mux);
and (n764, n740, n746);
xnor (n764_xnor, n764, n764);
or (n765_1, n763_mux, n764_mux);
or (n765, n762_mux, n765_1);
or (n765_1, n763, n764);
or (n765, n762, n765_1);
xnor (n765_xnor, n765, n765);
and (n782, n760_mux, n765_mux);
and (n782, n760, n765);
xnor (n782_xnor, n782, n782);
and (n783, n759_mux, n765_mux);
and (n783, n759, n765);
xnor (n783_xnor, n783, n783);
or (n784_1, n782_mux, n783_mux);
or (n784, n781_mux, n784_1);
or (n784_1, n782, n783);
or (n784, n781, n784_1);
xnor (n784_xnor, n784, n784);
and (n801, n779_mux, n784_mux);
and (n801, n779, n784);
xnor (n801_xnor, n801, n801);
and (n802, n778_mux, n784_mux);
and (n802, n778, n784);
xnor (n802_xnor, n802, n802);
or (n803_1, n801_mux, n802_mux);
or (n803, n800_mux, n803_1);
or (n803_1, n801, n802);
or (n803, n800, n803_1);
xnor (n803_xnor, n803, n803);
and (n820, n798_mux, n803_mux);
and (n820, n798, n803);
xnor (n820_xnor, n820, n820);
and (n821, n797_mux, n803_mux);
and (n821, n797, n803);
xnor (n821_xnor, n821, n821);
or (n822_1, n820_mux, n821_mux);
or (n822, n819_mux, n822_1);
or (n822_1, n820, n821);
or (n822, n819, n822_1);
xnor (n822_xnor, n822, n822);
and (n836, n817_mux, n822_mux);
and (n836, n817, n822);
xnor (n836_xnor, n836, n836);
and (n837, n816_mux, n822_mux);
and (n837, n816, n822);
xnor (n837_xnor, n837, n837);
or (n838_1, n836_mux, n837_mux);
or (n838, n835_mux, n838_1);
or (n838_1, n836, n837);
or (n838, n835, n838_1);
xnor (n838_xnor, n838, n838);
buf(n839, n838_mux);
buf(n839, n838);
xnor (n839_xnor, n839, n839);
and (n26, n25_mux, n839_mux);
and (n26, n25, n839);
xnor (n26_xnor, n26, n26);
buf(n825, g349_mux);
buf(n825, g349);
xnor (n825_xnor, n825, n825);
xnor (g8_xnor, g8, g8);
buf(g357, g8_mux);
buf(g357, g8);
xnor (g357_xnor, g357, g357);
buf(n826, g357_mux);
buf(n826, g357);
xnor (n826_xnor, n826, n826);
and (n840, n825_mux, n826_mux);
and (n840, n825, n826);
xnor (n840_xnor, n840, n840);
buf(n806, g350_mux);
buf(n806, g350);
xnor (n806_xnor, n806, n806);
buf(n807, n28_mux);
buf(n807, n28);
xnor (n807_xnor, n807, n807);
and (n828, n806_mux, n807_mux);
and (n828, n806, n807);
xnor (n828_xnor, n828, n828);
buf(n787, g351_mux);
buf(n787, g351);
xnor (n787_xnor, n787, n787);
buf(n788, n29_mux);
buf(n788, n29);
xnor (n788_xnor, n788, n788);
and (n809, n787_mux, n788_mux);
and (n809, n787, n788);
xnor (n809_xnor, n809, n809);
buf(n768, g352_mux);
buf(n768, g352);
xnor (n768_xnor, n768, n768);
buf(n769, n30_mux);
buf(n769, n30);
xnor (n769_xnor, n769, n769);
and (n790, n768_mux, n769_mux);
and (n790, n768, n769);
xnor (n790_xnor, n790, n790);
buf(n749, g353_mux);
buf(n749, g353);
xnor (n749_xnor, n749, n749);
buf(n750, n31_mux);
buf(n750, n31);
xnor (n750_xnor, n750, n750);
and (n771, n749_mux, n750_mux);
and (n771, n749, n750);
xnor (n771_xnor, n771, n771);
buf(n730, g354_mux);
buf(n730, g354);
xnor (n730_xnor, n730, n730);
buf(n731, n32_mux);
buf(n731, n32);
xnor (n731_xnor, n731, n731);
and (n752, n730_mux, n731_mux);
and (n752, n730, n731);
xnor (n752_xnor, n752, n752);
buf(n714, g355_mux);
buf(n714, g355);
xnor (n714_xnor, n714, n714);
buf(n715, n33_mux);
buf(n715, n33);
xnor (n715_xnor, n715, n715);
and (n733, n714_mux, n715_mux);
and (n733, n714, n715);
xnor (n733_xnor, n733, n733);
buf(n302, g356_mux);
buf(n302, g356);
xnor (n302_xnor, n302, n302);
buf(n303, n34_mux);
buf(n303, n34);
xnor (n303_xnor, n303, n303);
and (n717, n302_mux, n303_mux);
and (n717, n302, n303);
xnor (n717_xnor, n717, n717);
and (n734, n715_mux, n717_mux);
and (n734, n715, n717);
xnor (n734_xnor, n734, n734);
and (n735, n714_mux, n717_mux);
and (n735, n714, n717);
xnor (n735_xnor, n735, n735);
or (n736_1, n734_mux, n735_mux);
or (n736, n733_mux, n736_1);
or (n736_1, n734, n735);
or (n736, n733, n736_1);
xnor (n736_xnor, n736, n736);
and (n753, n731_mux, n736_mux);
and (n753, n731, n736);
xnor (n753_xnor, n753, n753);
and (n754, n730_mux, n736_mux);
and (n754, n730, n736);
xnor (n754_xnor, n754, n754);
or (n755_1, n753_mux, n754_mux);
or (n755, n752_mux, n755_1);
or (n755_1, n753, n754);
or (n755, n752, n755_1);
xnor (n755_xnor, n755, n755);
and (n772, n750_mux, n755_mux);
and (n772, n750, n755);
xnor (n772_xnor, n772, n772);
and (n773, n749_mux, n755_mux);
and (n773, n749, n755);
xnor (n773_xnor, n773, n773);
or (n774_1, n772_mux, n773_mux);
or (n774, n771_mux, n774_1);
or (n774_1, n772, n773);
or (n774, n771, n774_1);
xnor (n774_xnor, n774, n774);
and (n791, n769_mux, n774_mux);
and (n791, n769, n774);
xnor (n791_xnor, n791, n791);
and (n792, n768_mux, n774_mux);
and (n792, n768, n774);
xnor (n792_xnor, n792, n792);
or (n793_1, n791_mux, n792_mux);
or (n793, n790_mux, n793_1);
or (n793_1, n791, n792);
or (n793, n790, n793_1);
xnor (n793_xnor, n793, n793);
and (n810, n788_mux, n793_mux);
and (n810, n788, n793);
xnor (n810_xnor, n810, n810);
and (n811, n787_mux, n793_mux);
and (n811, n787, n793);
xnor (n811_xnor, n811, n811);
or (n812_1, n810_mux, n811_mux);
or (n812, n809_mux, n812_1);
or (n812_1, n810, n811);
or (n812, n809, n812_1);
xnor (n812_xnor, n812, n812);
and (n829, n807_mux, n812_mux);
and (n829, n807, n812);
xnor (n829_xnor, n829, n829);
and (n830, n806_mux, n812_mux);
and (n830, n806, n812);
xnor (n830_xnor, n830, n830);
or (n831_1, n829_mux, n830_mux);
or (n831, n828_mux, n831_1);
or (n831_1, n829, n830);
or (n831, n828, n831_1);
xnor (n831_xnor, n831, n831);
and (n841, n826_mux, n831_mux);
and (n841, n826, n831);
xnor (n841_xnor, n841, n841);
and (n842, n825_mux, n831_mux);
and (n842, n825, n831);
xnor (n842_xnor, n842, n842);
or (n843_1, n841_mux, n842_mux);
or (n843, n840_mux, n843_1);
or (n843_1, n841, n842);
or (n843, n840, n843_1);
xnor (n843_xnor, n843, n843);
buf(n844, n843_mux);
buf(n844, n843);
xnor (n844_xnor, n844, n844);
and (n27, n844_mux, n706_mux);
and (n27, n844, n706);
xnor (n27_xnor, n27, n27);
or (n845, n26_mux, n27_mux);
or (n845, n26, n27);
xnor (n845_xnor, n845, n845);
buf(n1454, n845_mux);
buf(n1454, n845);
xnor (n1454_xnor, n1454, n1454);
xor (n1346, n1315_mux, n1318_mux);
xor (n1346, n1315, n1318);
xnor (n1346_xnor, n1346, n1346);
buf(n1347, n1346_mux);
buf(n1347, n1346);
xnor (n1347_xnor, n1347, n1347);
buf(n1470, n1347_mux);
buf(n1470, n1347);
xnor (n1470_xnor, n1470, n1470);
and (n1478, n1454_mux, n1470_mux);
and (n1478, n1454, n1470);
xnor (n1478_xnor, n1478, n1478);
not(n22, n706_mux);
not(n22, n706);
xnor (n22_xnor, n22, n22);
xor (n818, n816_mux, n817_mux);
xor (n818, n816, n817);
xnor (n818_xnor, n818, n818);
xor (n823, n818_mux, n822_mux);
xor (n823, n818, n822);
xnor (n823_xnor, n823, n823);
buf(n824, n823_mux);
buf(n824, n823);
xnor (n824_xnor, n824, n824);
and (n23, n22_mux, n824_mux);
and (n23, n22, n824);
xnor (n23_xnor, n23, n23);
xor (n827, n825_mux, n826_mux);
xor (n827, n825, n826);
xnor (n827_xnor, n827, n827);
xor (n832, n827_mux, n831_mux);
xor (n832, n827, n831);
xnor (n832_xnor, n832, n832);
buf(n833, n832_mux);
buf(n833, n832);
xnor (n833_xnor, n833, n833);
and (n24, n833_mux, n706_mux);
and (n24, n833, n706);
xnor (n24_xnor, n24, n24);
or (n834, n23_mux, n24_mux);
or (n834, n23, n24);
xnor (n834_xnor, n834, n834);
buf(n1455, n834_mux);
buf(n1455, n834);
xnor (n1455_xnor, n1455, n1455);
and (n1479, n1455_mux, t_1);
and (n1479, n1455, t_1);
xnor (n1479_xnor, n1479, n1479);
not(n19, n706_mux);
not(n19, n706);
xnor (n19_xnor, n19, n19);
xor (n799, n797_mux, n798_mux);
xor (n799, n797, n798);
xnor (n799_xnor, n799, n799);
xor (n804, n799_mux, n803_mux);
xor (n804, n799, n803);
xnor (n804_xnor, n804, n804);
buf(n805, n804_mux);
buf(n805, n804);
xnor (n805_xnor, n805, n805);
and (n20, n19_mux, n805_mux);
and (n20, n19, n805);
xnor (n20_xnor, n20, n20);
xor (n808, n806_mux, n807_mux);
xor (n808, n806, n807);
xnor (n808_xnor, n808, n808);
xor (n813, n808_mux, n812_mux);
xor (n813, n808, n812);
xnor (n813_xnor, n813, n813);
buf(n814, n813_mux);
buf(n814, n813);
xnor (n814_xnor, n814, n814);
and (n21, n814_mux, n706_mux);
and (n21, n814, n706);
xnor (n21_xnor, n21, n21);
or (n815, n20_mux, n21_mux);
or (n815, n20, n21);
xnor (n815_xnor, n815, n815);
buf(n1456, n815_mux);
buf(n1456, n815);
xnor (n1456_xnor, n1456, n1456);
buf(n1471, n639_mux);
buf(n1471, n639);
xnor (n1471_xnor, n1471, n1471);
and (n1480, n1456_mux, n1471_mux);
and (n1480, n1456, n1471);
xnor (n1480_xnor, n1480, n1480);
not(n16, n706_mux);
not(n16, n706);
xnor (n16_xnor, n16, n16);
xor (n780, n778_mux, n779_mux);
xor (n780, n778, n779);
xnor (n780_xnor, n780, n780);
xor (n785, n780_mux, n784_mux);
xor (n785, n780, n784);
xnor (n785_xnor, n785, n785);
buf(n786, n785_mux);
buf(n786, n785);
xnor (n786_xnor, n786, n786);
and (n17, n16_mux, n786_mux);
and (n17, n16, n786);
xnor (n17_xnor, n17, n17);
xor (n789, n787_mux, n788_mux);
xor (n789, n787, n788);
xnor (n789_xnor, n789, n789);
xor (n794, n789_mux, n793_mux);
xor (n794, n789, n793);
xnor (n794_xnor, n794, n794);
buf(n795, n794_mux);
buf(n795, n794);
xnor (n795_xnor, n795, n795);
and (n18, n795_mux, n706_mux);
and (n18, n795, n706);
xnor (n18_xnor, n18, n18);
or (n796, n17_mux, n18_mux);
or (n796, n17, n18);
xnor (n796_xnor, n796, n796);
buf(n1457, n796_mux);
buf(n1457, n796);
xnor (n1457_xnor, n1457, n1457);
buf(n1472, n646_mux);
buf(n1472, n646);
xnor (n1472_xnor, n1472, n1472);
and (n1481, n1457_mux, n1472_mux);
and (n1481, n1457, n1472);
xnor (n1481_xnor, n1481, n1481);
not(n13, n706_mux);
not(n13, n706);
xnor (n13_xnor, n13, n13);
xor (n761, n759_mux, n760_mux);
xor (n761, n759, n760);
xnor (n761_xnor, n761, n761);
xor (n766, n761_mux, n765_mux);
xor (n766, n761, n765);
xnor (n766_xnor, n766, n766);
buf(n767, n766_mux);
buf(n767, n766);
xnor (n767_xnor, n767, n767);
and (n14, n13_mux, n767_mux);
and (n14, n13, n767);
xnor (n14_xnor, n14, n14);
xor (n770, n768_mux, n769_mux);
xor (n770, n768, n769);
xnor (n770_xnor, n770, n770);
xor (n775, n770_mux, n774_mux);
xor (n775, n770, n774);
xnor (n775_xnor, n775, n775);
buf(n776, n775_mux);
buf(n776, n775);
xnor (n776_xnor, n776, n776);
and (n15, n776_mux, n706_mux);
and (n15, n776, n706);
xnor (n15_xnor, n15, n15);
or (n777, n14_mux, n15_mux);
or (n777, n14, n15);
xnor (n777_xnor, n777, n777);
buf(n1458, n777_mux);
buf(n1458, n777);
xnor (n1458_xnor, n1458, n1458);
buf(n1473, n653_mux);
buf(n1473, n653);
xnor (n1473_xnor, n1473, n1473);
and (n1482, n1458_mux, n1473_mux);
and (n1482, n1458, n1473);
xnor (n1482_xnor, n1482, n1482);
not(n10, n706_mux);
not(n10, n706);
xnor (n10_xnor, n10, n10);
xor (n742, n740_mux, n741_mux);
xor (n742, n740, n741);
xnor (n742_xnor, n742, n742);
xor (n747, n742_mux, n746_mux);
xor (n747, n742, n746);
xnor (n747_xnor, n747, n747);
buf(n748, n747_mux);
buf(n748, n747);
xnor (n748_xnor, n748, n748);
and (n11, n10_mux, n748_mux);
and (n11, n10, n748);
xnor (n11_xnor, n11, n11);
xor (n751, n749_mux, n750_mux);
xor (n751, n749, n750);
xnor (n751_xnor, n751, n751);
xor (n756, n751_mux, n755_mux);
xor (n756, n751, n755);
xnor (n756_xnor, n756, n756);
buf(n757, n756_mux);
buf(n757, n756);
xnor (n757_xnor, n757, n757);
and (n12, n757_mux, n706_mux);
and (n12, n757, n706);
xnor (n12_xnor, n12, n12);
or (n758, n11_mux, n12_mux);
or (n758, n11, n12);
xnor (n758_xnor, n758, n758);
buf(n1459, n758_mux);
buf(n1459, n758);
xnor (n1459_xnor, n1459, n1459);
buf(n1474, n660_mux);
buf(n1474, n660);
xnor (n1474_xnor, n1474, n1474);
and (n1483, n1459_mux, n1474_mux);
and (n1483, n1459, n1474);
xnor (n1483_xnor, n1483, n1483);
not(n7, n706_mux);
not(n7, n706);
xnor (n7_xnor, n7, n7);
xor (n723, n721_mux, n722_mux);
xor (n723, n721, n722);
xnor (n723_xnor, n723, n723);
xor (n728, n723_mux, n727_mux);
xor (n728, n723, n727);
xnor (n728_xnor, n728, n728);
buf(n729, n728_mux);
buf(n729, n728);
xnor (n729_xnor, n729, n729);
and (n8, n7_mux, n729_mux);
and (n8, n7, n729);
xnor (n8_xnor, n8, n8);
xor (n732, n730_mux, n731_mux);
xor (n732, n730, n731);
xnor (n732_xnor, n732, n732);
xor (n737, n732_mux, n736_mux);
xor (n737, n732, n736);
xnor (n737_xnor, n737, n737);
buf(n738, n737_mux);
buf(n738, n737);
xnor (n738_xnor, n738, n738);
and (n9, n738_mux, n706_mux);
and (n9, n738, n706);
xnor (n9_xnor, n9, n9);
or (n739, n8_mux, n9_mux);
or (n739, n8, n9);
xnor (n739_xnor, n739, n739);
buf(n1460, n739_mux);
buf(n1460, n739);
xnor (n1460_xnor, n1460, n1460);
buf(n1475, n667_mux);
buf(n1475, n667);
xnor (n1475_xnor, n1475, n1475);
and (n1484, n1460_mux, n1475_mux);
and (n1484, n1460, n1475);
xnor (n1484_xnor, n1484, n1484);
not(n4, n706_mux);
not(n4, n706);
xnor (n4_xnor, n4, n4);
xor (n710, n708_mux, n709_mux);
xor (n710, n708, n709);
xnor (n710_xnor, n710, n710);
xor (n712, n710_mux, n711_mux);
xor (n712, n710, n711);
xnor (n712_xnor, n712, n712);
buf(n713, n712_mux);
buf(n713, n712);
xnor (n713_xnor, n713, n713);
and (n5, n4_mux, n713_mux);
and (n5, n4, n713);
xnor (n5_xnor, n5, n5);
xor (n716, n714_mux, n715_mux);
xor (n716, n714, n715);
xnor (n716_xnor, n716, n716);
xor (n718, n716_mux, n717_mux);
xor (n718, n716, n717);
xnor (n718_xnor, n718, n718);
buf(n719, n718_mux);
buf(n719, n718);
xnor (n719_xnor, n719, n719);
and (n6, n719_mux, n706_mux);
and (n6, n719, n706);
xnor (n6_xnor, n6, n6);
or (n720, n5_mux, n6_mux);
or (n720, n5, n6);
xnor (n720_xnor, n720, n720);
buf(n1461, n720_mux);
buf(n1461, n720);
xnor (n1461_xnor, n1461, n1461);
buf(n1476, n674_mux);
buf(n1476, n674);
xnor (n1476_xnor, n1476, n1476);
and (n1485, n1461_mux, n1476_mux);
and (n1485, n1461, n1476);
xnor (n1485_xnor, n1485, n1485);
not(n1, n706_mux);
not(n1, n706);
xnor (n1_xnor, n1, n1);
xor (n300, n298_mux, n299_mux);
xor (n300, n298, n299);
xnor (n300_xnor, n300, n300);
buf(n301, n300_mux);
buf(n301, n300);
xnor (n301_xnor, n301, n301);
and (n2, n1_mux, n301_mux);
and (n2, n1, n301);
xnor (n2_xnor, n2, n2);
xor (n304, n302_mux, n303_mux);
xor (n304, n302, n303);
xnor (n304_xnor, n304, n304);
buf(n305, n304_mux);
buf(n305, n304);
xnor (n305_xnor, n305, n305);
and (n3, n305_mux, n706_mux);
and (n3, n305, n706);
xnor (n3_xnor, n3, n3);
or (n707, n2_mux, n3_mux);
or (n707, n2, n3);
xnor (n707_xnor, n707, n707);
buf(n1462, n707_mux);
buf(n1462, n707);
xnor (n1462_xnor, n1462, n1462);
buf(n1477, n681_mux);
buf(n1477, n681);
xnor (n1477_xnor, n1477, n1477);
and (n1486, n1462_mux, n1477_mux);
and (n1486, n1462, n1477);
xnor (n1486_xnor, n1486, n1486);
and (n1487, n1476_mux, n1486_mux);
and (n1487, n1476, n1486);
xnor (n1487_xnor, n1487, n1487);
and (n1488, n1461_mux, n1486_mux);
and (n1488, n1461, n1486);
xnor (n1488_xnor, n1488, n1488);
or (n1489_1, n1487_mux, n1488_mux);
or (n1489, n1485_mux, n1489_1);
or (n1489_1, n1487, n1488);
or (n1489, n1485, n1489_1);
xnor (n1489_xnor, n1489, n1489);
and (n1490, n1475_mux, n1489_mux);
and (n1490, n1475, n1489);
xnor (n1490_xnor, n1490, n1490);
and (n1491, n1460_mux, n1489_mux);
and (n1491, n1460, n1489);
xnor (n1491_xnor, n1491, n1491);
or (n1492_1, n1490_mux, n1491_mux);
or (n1492, n1484_mux, n1492_1);
or (n1492_1, n1490, n1491);
or (n1492, n1484, n1492_1);
xnor (n1492_xnor, n1492, n1492);
and (n1493, n1474_mux, n1492_mux);
and (n1493, n1474, n1492);
xnor (n1493_xnor, n1493, n1493);
and (n1494, n1459_mux, n1492_mux);
and (n1494, n1459, n1492);
xnor (n1494_xnor, n1494, n1494);
or (n1495_1, n1493_mux, n1494_mux);
or (n1495, n1483_mux, n1495_1);
or (n1495_1, n1493, n1494);
or (n1495, n1483, n1495_1);
xnor (n1495_xnor, n1495, n1495);
and (n1496, n1473_mux, n1495_mux);
and (n1496, n1473, n1495);
xnor (n1496_xnor, n1496, n1496);
and (n1497, n1458_mux, n1495_mux);
and (n1497, n1458, n1495);
xnor (n1497_xnor, n1497, n1497);
or (n1498_1, n1496_mux, n1497_mux);
or (n1498, n1482_mux, n1498_1);
or (n1498_1, n1496, n1497);
or (n1498, n1482, n1498_1);
xnor (n1498_xnor, n1498, n1498);
and (n1499, n1472_mux, n1498_mux);
and (n1499, n1472, n1498);
xnor (n1499_xnor, n1499, n1499);
and (n1500, n1457_mux, n1498_mux);
and (n1500, n1457, n1498);
xnor (n1500_xnor, n1500, n1500);
or (n1501_1, n1499_mux, n1500_mux);
or (n1501, n1481_mux, n1501_1);
or (n1501_1, n1499, n1500);
or (n1501, n1481, n1501_1);
xnor (n1501_xnor, n1501, n1501);
and (n1502, n1471_mux, n1501_mux);
and (n1502, n1471, n1501);
xnor (n1502_xnor, n1502, n1502);
and (n1503, n1456_mux, n1501_mux);
and (n1503, n1456, n1501);
xnor (n1503_xnor, n1503, n1503);
or (n1504_1, n1502_mux, n1503_mux);
or (n1504, n1480_mux, n1504_1);
or (n1504_1, n1502, n1503);
or (n1504, n1480, n1504_1);
xnor (n1504_xnor, n1504, n1504);
and (n1505, t_1, n1504_mux);
and (n1505, t_1, n1504);
xnor (n1505_xnor, n1505, n1505);
and (n1506, n1455_mux, n1504_mux);
and (n1506, n1455, n1504);
xnor (n1506_xnor, n1506, n1506);
or (n1507_1, n1505_mux, n1506_mux);
or (n1507, n1479_mux, n1507_1);
or (n1507_1, n1505, n1506);
or (n1507, n1479, n1507_1);
xnor (n1507_xnor, n1507, n1507);
and (n1508, n1470_mux, n1507_mux);
and (n1508, n1470, n1507);
xnor (n1508_xnor, n1508, n1508);
and (n1509, n1454_mux, n1507_mux);
and (n1509, n1454, n1507);
xnor (n1509_xnor, n1509, n1509);
or (n1510_1, n1508_mux, n1509_mux);
or (n1510, n1478_mux, n1510_1);
or (n1510_1, n1508, n1509);
or (n1510, n1478, n1510_1);
xnor (n1510_xnor, n1510, n1510);
and (n1511, n1469_mux, n1510_mux);
and (n1511, n1469, n1510);
xnor (n1511_xnor, n1511, n1511);
and (n1512, n1468_mux, n1511_mux);
and (n1512, n1468, n1511);
xnor (n1512_xnor, n1512, n1512);
and (n1513, n1467_mux, n1512_mux);
and (n1513, n1467, n1512);
xnor (n1513_xnor, n1513, n1513);
and (n1514, n1466_mux, n1513_mux);
and (n1514, n1466, n1513);
xnor (n1514_xnor, n1514, n1514);
and (n1515, n1465_mux, n1514_mux);
and (n1515, n1465, n1514);
xnor (n1515_xnor, n1515, n1515);
and (n1516, n1464_mux, n1515_mux);
and (n1516, n1464, n1515);
xnor (n1516_xnor, n1516, n1516);
and (n1517, n1463_mux, n1516_mux);
and (n1517, n1463, n1516);
xnor (n1517_xnor, n1517, n1517);
buf(n1518, n1517_mux);
buf(n1518, n1517);
xnor (n1518_xnor, n1518, n1518);
buf(n99, n1518_mux);
buf(g80, n99);
buf(n99, n1518);
buf(g80, n99);
xnor (g80_xnor, g80, g80);
xor (n1519, n1463_mux, n1516_mux);
xor (n1519, n1463, n1516);
xnor (n1519_xnor, n1519, n1519);
buf(n1520, n1519_mux);
buf(n1520, n1519);
xnor (n1520_xnor, n1520, n1520);
buf(n100, n1520_mux);
buf(g81, n100);
buf(n100, n1520);
buf(g81, n100);
xnor (g81_xnor, g81, g81);
xor (n1521, n1464_mux, n1515_mux);
xor (n1521, n1464, n1515);
xnor (n1521_xnor, n1521, n1521);
buf(n1522, n1521_mux);
buf(n1522, n1521);
xnor (n1522_xnor, n1522, n1522);
buf(n101, n1522_mux);
buf(g82, n101);
buf(n101, n1522);
buf(g82, n101);
xnor (g82_xnor, g82, g82);
xor (n1523, n1465_mux, n1514_mux);
xor (n1523, n1465, n1514);
xnor (n1523_xnor, n1523, n1523);
buf(n1524, n1523_mux);
buf(n1524, n1523);
xnor (n1524_xnor, n1524, n1524);
buf(n102, n1524_mux);
buf(g83, n102);
buf(n102, n1524);
buf(g83, n102);
xnor (g83_xnor, g83, g83);
xor (n1525, n1466_mux, n1513_mux);
xor (n1525, n1466, n1513);
xnor (n1525_xnor, n1525, n1525);
buf(n1526, n1525_mux);
buf(n1526, n1525);
xnor (n1526_xnor, n1526, n1526);
buf(n103, n1526_mux);
buf(g84, n103);
buf(n103, n1526);
buf(g84, n103);
xnor (g84_xnor, g84, g84);
xor (n1527, n1467_mux, n1512_mux);
xor (n1527, n1467, n1512);
xnor (n1527_xnor, n1527, n1527);
buf(n1528, n1527_mux);
buf(n1528, n1527);
xnor (n1528_xnor, n1528, n1528);
buf(n104, n1528_mux);
buf(g85, n104);
buf(n104, n1528);
buf(g85, n104);
xnor (g85_xnor, g85, g85);
xor (n1529, n1468_mux, n1511_mux);
xor (n1529, n1468, n1511);
xnor (n1529_xnor, n1529, n1529);
buf(n1530, n1529_mux);
buf(n1530, n1529);
xnor (n1530_xnor, n1530, n1530);
buf(n105, n1530_mux);
buf(g86, n105);
buf(n105, n1530);
buf(g86, n105);
xnor (g86_xnor, g86, g86);
xor (n1531, n1469_mux, n1510_mux);
xor (n1531, n1469, n1510);
xnor (n1531_xnor, n1531, n1531);
buf(n1532, n1531_mux);
buf(n1532, n1531);
xnor (n1532_xnor, n1532, n1532);
buf(n106, n1532_mux);
buf(g87, n106);
buf(n106, n1532);
buf(g87, n106);
xnor (g87_xnor, g87, g87);
xor (n1533, n1454_mux, n1470_mux);
xor (n1533, n1454, n1470);
xnor (n1533_xnor, n1533, n1533);
xor (n1534, n1533_mux, n1507_mux);
xor (n1534, n1533, n1507);
xnor (n1534_xnor, n1534, n1534);
buf(n1535, n1534_mux);
buf(n1535, n1534);
xnor (n1535_xnor, n1535, n1535);
buf(n107, n1535_mux);
buf(g88, n107);
buf(n107, n1535);
buf(g88, n107);
xnor (g88_xnor, g88, g88);
xor (n1536, n1455_mux, t_1);
xor (n1536, n1455, t_1);
xnor (n1536_xnor, n1536, n1536);
xor (n1537, n1536_mux, n1504_mux);
xor (n1537, n1536, n1504);
xnor (n1537_xnor, n1537, n1537);
buf(n1538, n1537_mux);
buf(n1538, n1537);
xnor (n1538_xnor, n1538, n1538);
buf(n108, n1538_mux);
buf(g89, n108);
buf(n108, n1538);
buf(g89, n108);
xnor (g89_xnor, g89, g89);
xor (n1539, n1456_mux, n1471_mux);
xor (n1539, n1456, n1471);
xnor (n1539_xnor, n1539, n1539);
xor (n1540, n1539_mux, n1501_mux);
xor (n1540, n1539, n1501);
xnor (n1540_xnor, n1540, n1540);
buf(n1541, n1540_mux);
buf(n1541, n1540);
xnor (n1541_xnor, n1541, n1541);
buf(n109, n1541_mux);
buf(g90, n109);
buf(n109, n1541);
buf(g90, n109);
xnor (g90_xnor, g90, g90);
xor (n1542, n1457_mux, n1472_mux);
xor (n1542, n1457, n1472);
xnor (n1542_xnor, n1542, n1542);
xor (n1543, n1542_mux, n1498_mux);
xor (n1543, n1542, n1498);
xnor (n1543_xnor, n1543, n1543);
buf(n1544, n1543_mux);
buf(n1544, n1543);
xnor (n1544_xnor, n1544, n1544);
buf(n110, n1544_mux);
buf(g91, n110);
buf(n110, n1544);
buf(g91, n110);
xnor (g91_xnor, g91, g91);
xor (n1545, n1458_mux, n1473_mux);
xor (n1545, n1458, n1473);
xnor (n1545_xnor, n1545, n1545);
xor (n1546, n1545_mux, n1495_mux);
xor (n1546, n1545, n1495);
xnor (n1546_xnor, n1546, n1546);
buf(n1547, n1546_mux);
buf(n1547, n1546);
xnor (n1547_xnor, n1547, n1547);
buf(n111, n1547_mux);
buf(g92, n111);
buf(n111, n1547);
buf(g92, n111);
xnor (g92_xnor, g92, g92);
xor (n1548, n1459_mux, n1474_mux);
xor (n1548, n1459, n1474);
xnor (n1548_xnor, n1548, n1548);
xor (n1549, n1548_mux, n1492_mux);
xor (n1549, n1548, n1492);
xnor (n1549_xnor, n1549, n1549);
buf(n1550, n1549_mux);
buf(n1550, n1549);
xnor (n1550_xnor, n1550, n1550);
buf(n112, n1550_mux);
buf(g93, n112);
buf(n112, n1550);
buf(g93, n112);
xnor (g93_xnor, g93, g93);
xor (n1551, n1460_mux, n1475_mux);
xor (n1551, n1460, n1475);
xnor (n1551_xnor, n1551, n1551);
xor (n1552, n1551_mux, n1489_mux);
xor (n1552, n1551, n1489);
xnor (n1552_xnor, n1552, n1552);
buf(n1553, n1552_mux);
buf(n1553, n1552);
xnor (n1553_xnor, n1553, n1553);
buf(n113, n1553_mux);
buf(g94, n113);
buf(n113, n1553);
buf(g94, n113);
xnor (g94_xnor, g94, g94);
xor (n1554, n1461_mux, n1476_mux);
xor (n1554, n1461, n1476);
xnor (n1554_xnor, n1554, n1554);
xor (n1555, n1554_mux, n1486_mux);
xor (n1555, n1554, n1486);
xnor (n1555_xnor, n1555, n1555);
buf(n1556, n1555_mux);
buf(n1556, n1555);
xnor (n1556_xnor, n1556, n1556);
buf(n114, n1556_mux);
buf(g95, n114);
buf(n114, n1556);
buf(g95, n114);
xnor (g95_xnor, g95, g95);
xor (n1557, n1462_mux, n1477_mux);
xor (n1557, n1462, n1477);
xnor (n1557_xnor, n1557, n1557);
buf(n1558, n1557_mux);
buf(n1558, n1557);
xnor (n1558_xnor, n1558, n1558);
buf(n115, n1558_mux);
buf(g96, n115);
buf(n115, n1558);
buf(g96, n115);
xnor (g96_xnor, g96, g96);
buf(n116, 1'b0);
buf(g97, n116);
buf(n117, 1'b0);
buf(g98, n117);
buf(n118, 1'b0);
buf(g99, n118);
buf(n119, 1'b0);
buf(g100, n119);
buf(n120, 1'b0);
buf(g101, n120);
buf(n121, 1'b0);
buf(g102, n121);
buf(n122, 1'b0);
buf(g103, n122);
buf(n123, 1'b0);
buf(g104, n123);
buf(n124, 1'b0);
buf(g105, n124);
buf(n125, 1'b0);
buf(g106, n125);
buf(n126, 1'b0);
buf(g107, n126);
buf(n127, 1'b0);
buf(g108, n127);
buf(n128, 1'b0);
buf(g109, n128);
buf(n129, 1'b0);
buf(g110, n129);
buf(n130, 1'b0);
buf(g111, n130);
buf(n131, 1'b0);
buf(g112, n131);
buf(n132, 1'b0);
buf(g113, n132);
buf(n133, 1'b0);
buf(g114, n133);
buf(n134, 1'b0);
buf(g115, n134);
buf(n135, 1'b0);
buf(g116, n135);
buf(n136, 1'b0);
buf(g117, n136);
buf(n137, 1'b0);
buf(g118, n137);
buf(n138, 1'b0);
buf(g119, n138);
buf(n139, 1'b0);
buf(g120, n139);
buf(n140, 1'b0);
buf(g121, n140);
buf(n141, 1'b0);
buf(g122, n141);
buf(n142, 1'b0);
buf(g123, n142);
buf(n143, 1'b0);
buf(g124, n143);
buf(n144, 1'b0);
buf(g125, n144);
buf(n145, 1'b0);
buf(g126, n145);
buf(n146, 1'b0);
buf(g127, n146);
buf(n147, 1'b0);
buf(g128, n147);
buf(n148, 1'b0);
buf(g129, n148);
buf(n149, 1'b0);
buf(g130, n149);
buf(n150, 1'b0);
buf(g131, n150);
buf(n151, 1'b0);
buf(g132, n151);
buf(n152, 1'b0);
buf(g133, n152);
buf(n153, 1'b0);
buf(g134, n153);
buf(n154, 1'b0);
buf(g135, n154);
buf(n155, 1'b0);
buf(g136, n155);
buf(n156, 1'b0);
buf(g137, n156);
buf(n157, 1'b0);
buf(g138, n157);
buf(n158, 1'b0);
buf(g139, n158);
buf(n159, 1'b0);
buf(g140, n159);
buf(n160, 1'b0);
buf(g141, n160);
buf(n161, 1'b0);
buf(g142, n161);
buf(n162, 1'b0);
buf(g143, n162);
buf(n549, g357_mux);
buf(n549, g357);
xnor (n549_xnor, n549, n549);
buf(n545, n43_mux);
buf(n545, n43);
xnor (n545_xnor, n545, n545);
and (n866, n549_mux, n545_mux);
and (n866, n549, n545);
xnor (n866_xnor, n866, n866);
not(n867, n490_mux);
not(n867, n490);
xnor (n867_xnor, n867, n867);
not(n546, n545_mux);
not(n546, n545);
xnor (n546_xnor, n546, n546);
and (n868, n546_mux, n490_mux);
and (n868, n546, n490);
xnor (n868_xnor, n868, n868);
nor (n869, n867_mux, n868_mux);
nor (n869, n867, n868);
xnor (n869_xnor, n869, n869);
and (n870, n499_mux, n472_mux);
and (n870, n499, n472);
xnor (n870_xnor, n870, n870);
and (n871, n869_mux, n870_mux);
and (n871, n869, n870);
xnor (n871_xnor, n871, n871);
and (n872, n515_mux, n475_mux);
and (n872, n515, n475);
xnor (n872_xnor, n872, n872);
and (n873, n870_mux, n872_mux);
and (n873, n870, n872);
xnor (n873_xnor, n873, n873);
and (n874, n869_mux, n872_mux);
and (n874, n869, n872);
xnor (n874_xnor, n874, n874);
or (n875_1, n873_mux, n874_mux);
or (n875, n871_mux, n875_1);
or (n875_1, n873, n874);
or (n875, n871, n875_1);
xnor (n875_xnor, n875, n875);
not(n876, n499_mux);
not(n876, n499);
xnor (n876_xnor, n876, n876);
and (n877, n546_mux, n499_mux);
and (n877, n546, n499);
xnor (n877_xnor, n877, n877);
nor (n878, n876_mux, n877_mux);
nor (n878, n876, n877);
xnor (n878_xnor, n878, n878);
and (n879, n875_mux, n878_mux);
and (n879, n875, n878);
xnor (n879_xnor, n879, n879);
and (n880, n515_mux, n472_mux);
and (n880, n515, n472);
xnor (n880_xnor, n880, n880);
and (n881, n878_mux, n880_mux);
and (n881, n878, n880);
xnor (n881_xnor, n881, n881);
and (n882, n875_mux, n880_mux);
and (n882, n875, n880);
xnor (n882_xnor, n882, n882);
or (n883_1, n881_mux, n882_mux);
or (n883, n879_mux, n883_1);
or (n883_1, n881, n882);
or (n883, n879, n883_1);
xnor (n883_xnor, n883, n883);
not(n884, n515_mux);
not(n884, n515);
xnor (n884_xnor, n884, n884);
and (n885, n546_mux, n515_mux);
and (n885, n546, n515);
xnor (n885_xnor, n885, n885);
nor (n886, n884_mux, n885_mux);
nor (n886, n884, n885);
xnor (n886_xnor, n886, n886);
and (n887, n883_mux, n886_mux);
and (n887, n883, n886);
xnor (n887_xnor, n887, n887);
not(n550, n549_mux);
not(n550, n549);
xnor (n550_xnor, n550, n550);
and (n888, n550_mux, n472_mux);
and (n888, n550, n472);
xnor (n888_xnor, n888, n888);
not(n889, n472_mux);
not(n889, n472);
xnor (n889_xnor, n889, n889);
nor (n890, n888_mux, n889_mux);
nor (n890, n888, n889);
xnor (n890_xnor, n890, n890);
and (n891, n886_mux, n890_mux);
and (n891, n886, n890);
xnor (n891_xnor, n891, n891);
and (n892, n883_mux, n890_mux);
and (n892, n883, n890);
xnor (n892_xnor, n892, n892);
or (n893_1, n891_mux, n892_mux);
or (n893, n887_mux, n893_1);
or (n893_1, n891, n892);
or (n893, n887, n893_1);
xnor (n893_xnor, n893, n893);
and (n894, n866_mux, n893_mux);
and (n894, n866, n893);
xnor (n894_xnor, n894, n894);
xor (n895, n866_mux, n893_mux);
xor (n895, n866, n893);
xnor (n895_xnor, n895, n895);
xor (n896, n883_mux, n886_mux);
xor (n896, n883, n886);
xnor (n896_xnor, n896, n896);
xor (n897, n896_mux, n890_mux);
xor (n897, n896, n890);
xnor (n897_xnor, n897, n897);
not(n898, n486_mux);
not(n898, n486);
xnor (n898_xnor, n898, n898);
and (n899, n546_mux, n486_mux);
and (n899, n546, n486);
xnor (n899_xnor, n899, n899);
nor (n900, n898_mux, n899_mux);
nor (n900, n898, n899);
xnor (n900_xnor, n900, n900);
and (n901, n490_mux, n472_mux);
and (n901, n490, n472);
xnor (n901_xnor, n901, n901);
and (n902, n900_mux, n901_mux);
and (n902, n900, n901);
xnor (n902_xnor, n902, n902);
and (n903, n550_mux, n509_mux);
and (n903, n550, n509);
xnor (n903_xnor, n903, n903);
not(n904, n509_mux);
not(n904, n509);
xnor (n904_xnor, n904, n904);
nor (n905, n903_mux, n904_mux);
nor (n905, n903, n904);
xnor (n905_xnor, n905, n905);
and (n906, n901_mux, n905_mux);
and (n906, n901, n905);
xnor (n906_xnor, n906, n906);
and (n907, n900_mux, n905_mux);
and (n907, n900, n905);
xnor (n907_xnor, n907, n907);
or (n908_1, n906_mux, n907_mux);
or (n908, n902_mux, n908_1);
or (n908_1, n906, n907);
or (n908, n902, n908_1);
xnor (n908_xnor, n908, n908);
and (n909, n490_mux, n475_mux);
and (n909, n490, n475);
xnor (n909_xnor, n909, n909);
and (n910, n499_mux, n479_mux);
and (n910, n499, n479);
xnor (n910_xnor, n910, n910);
and (n911, n909_mux, n910_mux);
and (n911, n909, n910);
xnor (n911_xnor, n911, n911);
and (n912, n515_mux, n509_mux);
and (n912, n515, n509);
xnor (n912_xnor, n912, n912);
and (n913, n910_mux, n912_mux);
and (n913, n910, n912);
xnor (n913_xnor, n913, n913);
and (n914, n909_mux, n912_mux);
and (n914, n909, n912);
xnor (n914_xnor, n914, n914);
or (n915_1, n913_mux, n914_mux);
or (n915, n911_mux, n915_1);
or (n915_1, n913, n914);
or (n915, n911, n915_1);
xnor (n915_xnor, n915, n915);
and (n916, n499_mux, n475_mux);
and (n916, n499, n475);
xnor (n916_xnor, n916, n916);
and (n917, n915_mux, n916_mux);
and (n917, n915, n916);
xnor (n917_xnor, n917, n917);
and (n918, n515_mux, n479_mux);
and (n918, n515, n479);
xnor (n918_xnor, n918, n918);
and (n919, n916_mux, n918_mux);
and (n919, n916, n918);
xnor (n919_xnor, n919, n919);
and (n920, n915_mux, n918_mux);
and (n920, n915, n918);
xnor (n920_xnor, n920, n920);
or (n921_1, n919_mux, n920_mux);
or (n921, n917_mux, n921_1);
or (n921_1, n919, n920);
or (n921, n917, n921_1);
xnor (n921_xnor, n921, n921);
and (n922, n908_mux, n921_mux);
and (n922, n908, n921);
xnor (n922_xnor, n922, n922);
xor (n923, n869_mux, n870_mux);
xor (n923, n869, n870);
xnor (n923_xnor, n923, n923);
xor (n924, n923_mux, n872_mux);
xor (n924, n923, n872);
xnor (n924_xnor, n924, n924);
and (n925, n921_mux, n924_mux);
and (n925, n921, n924);
xnor (n925_xnor, n925, n925);
and (n926, n908_mux, n924_mux);
and (n926, n908, n924);
xnor (n926_xnor, n926, n926);
or (n927_1, n925_mux, n926_mux);
or (n927, n922_mux, n927_1);
or (n927_1, n925, n926);
or (n927, n922, n927_1);
xnor (n927_xnor, n927, n927);
and (n928, n550_mux, n475_mux);
and (n928, n550, n475);
xnor (n928_xnor, n928, n928);
not(n929, n475_mux);
not(n929, n475);
xnor (n929_xnor, n929, n929);
nor (n930, n928_mux, n929_mux);
nor (n930, n928, n929);
xnor (n930_xnor, n930, n930);
and (n931, n927_mux, n930_mux);
and (n931, n927, n930);
xnor (n931_xnor, n931, n931);
xor (n932, n875_mux, n878_mux);
xor (n932, n875, n878);
xnor (n932_xnor, n932, n932);
xor (n933, n932_mux, n880_mux);
xor (n933, n932, n880);
xnor (n933_xnor, n933, n933);
and (n934, n930_mux, n933_mux);
and (n934, n930, n933);
xnor (n934_xnor, n934, n934);
and (n935, n927_mux, n933_mux);
and (n935, n927, n933);
xnor (n935_xnor, n935, n935);
or (n936_1, n934_mux, n935_mux);
or (n936, n931_mux, n936_1);
or (n936_1, n934, n935);
or (n936, n931, n936_1);
xnor (n936_xnor, n936, n936);
and (n937, n897_mux, n936_mux);
and (n937, n897, n936);
xnor (n937_xnor, n937, n937);
xor (n938, n897_mux, n936_mux);
xor (n938, n897, n936);
xnor (n938_xnor, n938, n938);
xor (n939, n927_mux, n930_mux);
xor (n939, n927, n930);
xnor (n939_xnor, n939, n939);
xor (n940, n939_mux, n933_mux);
xor (n940, n939, n933);
xnor (n940_xnor, n940, n940);
and (n941, n490_mux, n479_mux);
and (n941, n490, n479);
xnor (n941_xnor, n941, n941);
and (n942, n499_mux, n509_mux);
and (n942, n499, n509);
xnor (n942_xnor, n942, n942);
and (n943, n941_mux, n942_mux);
and (n943, n941, n942);
xnor (n943_xnor, n943, n943);
and (n944, n515_mux, n484_mux);
and (n944, n515, n484);
xnor (n944_xnor, n944, n944);
and (n945, n942_mux, n944_mux);
and (n945, n942, n944);
xnor (n945_xnor, n945, n945);
and (n946, n941_mux, n944_mux);
and (n946, n941, n944);
xnor (n946_xnor, n946, n946);
or (n947_1, n945_mux, n946_mux);
or (n947, n943_mux, n947_1);
or (n947_1, n945, n946);
or (n947, n943, n947_1);
xnor (n947_xnor, n947, n947);
and (n948, n478_mux, n472_mux);
and (n948, n478, n472);
xnor (n948_xnor, n948, n948);
and (n949, n486_mux, n475_mux);
and (n949, n486, n475);
xnor (n949_xnor, n949, n949);
and (n950, n948_mux, n949_mux);
and (n950, n948, n949);
xnor (n950_xnor, n950, n950);
and (n951, n947_mux, n950_mux);
and (n951, n947, n950);
xnor (n951_xnor, n951, n951);
xor (n952, n909_mux, n910_mux);
xor (n952, n909, n910);
xnor (n952_xnor, n952, n952);
xor (n953, n952_mux, n912_mux);
xor (n953, n952, n912);
xnor (n953_xnor, n953, n953);
and (n954, n950_mux, n953_mux);
and (n954, n950, n953);
xnor (n954_xnor, n954, n954);
and (n955, n947_mux, n953_mux);
and (n955, n947, n953);
xnor (n955_xnor, n955, n955);
or (n956_1, n954_mux, n955_mux);
or (n956, n951_mux, n956_1);
or (n956_1, n954, n955);
or (n956, n951, n956_1);
xnor (n956_xnor, n956, n956);
xor (n957, n900_mux, n901_mux);
xor (n957, n900, n901);
xnor (n957_xnor, n957, n957);
xor (n958, n957_mux, n905_mux);
xor (n958, n957, n905);
xnor (n958_xnor, n958, n958);
and (n959, n956_mux, n958_mux);
and (n959, n956, n958);
xnor (n959_xnor, n959, n959);
xor (n960, n915_mux, n916_mux);
xor (n960, n915, n916);
xnor (n960_xnor, n960, n960);
xor (n961, n960_mux, n918_mux);
xor (n961, n960, n918);
xnor (n961_xnor, n961, n961);
and (n962, n958_mux, n961_mux);
and (n962, n958, n961);
xnor (n962_xnor, n962, n962);
and (n963, n956_mux, n961_mux);
and (n963, n956, n961);
xnor (n963_xnor, n963, n963);
or (n964_1, n962_mux, n963_mux);
or (n964, n959_mux, n964_1);
or (n964_1, n962, n963);
or (n964, n959, n964_1);
xnor (n964_xnor, n964, n964);
and (n965, n550_mux, n479_mux);
and (n965, n550, n479);
xnor (n965_xnor, n965, n965);
not(n966, n479_mux);
not(n966, n479);
xnor (n966_xnor, n966, n966);
nor (n967, n965_mux, n966_mux);
nor (n967, n965, n966);
xnor (n967_xnor, n967, n967);
and (n968, n964_mux, n967_mux);
and (n968, n964, n967);
xnor (n968_xnor, n968, n968);
xor (n969, n908_mux, n921_mux);
xor (n969, n908, n921);
xnor (n969_xnor, n969, n969);
xor (n970, n969_mux, n924_mux);
xor (n970, n969, n924);
xnor (n970_xnor, n970, n970);
and (n971, n967_mux, n970_mux);
and (n971, n967, n970);
xnor (n971_xnor, n971, n971);
and (n972, n964_mux, n970_mux);
and (n972, n964, n970);
xnor (n972_xnor, n972, n972);
or (n973_1, n971_mux, n972_mux);
or (n973, n968_mux, n973_1);
or (n973_1, n971, n972);
or (n973, n968, n973_1);
xnor (n973_xnor, n973, n973);
and (n974, n940_mux, n973_mux);
and (n974, n940, n973);
xnor (n974_xnor, n974, n974);
xor (n975, n940_mux, n973_mux);
xor (n975, n940, n973);
xnor (n975_xnor, n975, n975);
xor (n976, n964_mux, n967_mux);
xor (n976, n964, n967);
xnor (n976_xnor, n976, n976);
xor (n977, n976_mux, n970_mux);
xor (n977, n976, n970);
xnor (n977_xnor, n977, n977);
not(n978, n478_mux);
not(n978, n478);
xnor (n978_xnor, n978, n978);
and (n979, n546_mux, n478_mux);
and (n979, n546, n478);
xnor (n979_xnor, n979, n979);
nor (n980, n978_mux, n979_mux);
nor (n980, n978, n979);
xnor (n980_xnor, n980, n980);
and (n981, n486_mux, n472_mux);
and (n981, n486, n472);
xnor (n981_xnor, n981, n981);
and (n982, n980_mux, n981_mux);
and (n982, n980, n981);
xnor (n982_xnor, n982, n982);
and (n983, n550_mux, n484_mux);
and (n983, n550, n484);
xnor (n983_xnor, n983, n983);
not(n984, n484_mux);
not(n984, n484);
xnor (n984_xnor, n984, n984);
nor (n985, n983_mux, n984_mux);
nor (n985, n983, n984);
xnor (n985_xnor, n985, n985);
and (n986, n981_mux, n985_mux);
and (n986, n981, n985);
xnor (n986_xnor, n986, n986);
and (n987, n980_mux, n985_mux);
and (n987, n980, n985);
xnor (n987_xnor, n987, n987);
or (n988_1, n986_mux, n987_mux);
or (n988, n982_mux, n988_1);
or (n988_1, n986, n987);
or (n988, n982, n988_1);
xnor (n988_xnor, n988, n988);
and (n537, n490_mux, n509_mux);
and (n537, n490, n509);
xnor (n537_xnor, n537, n537);
and (n538, n499_mux, n484_mux);
and (n538, n499, n484);
xnor (n538_xnor, n538, n538);
and (n989, n537_mux, n538_mux);
and (n989, n537, n538);
xnor (n989_xnor, n989, n989);
and (n540, n515_mux, n487_mux);
and (n540, n515, n487);
xnor (n540_xnor, n540, n540);
and (n990, n538_mux, n540_mux);
and (n990, n538, n540);
xnor (n990_xnor, n990, n990);
and (n991, n537_mux, n540_mux);
and (n991, n537, n540);
xnor (n991_xnor, n991, n991);
or (n992_1, n990_mux, n991_mux);
or (n992, n989_mux, n992_1);
or (n992_1, n990, n991);
or (n992, n989, n992_1);
xnor (n992_xnor, n992, n992);
xor (n993, n941_mux, n942_mux);
xor (n993, n941, n942);
xnor (n993_xnor, n993, n993);
xor (n994, n993_mux, n944_mux);
xor (n994, n993, n944);
xnor (n994_xnor, n994, n994);
and (n995, n992_mux, n994_mux);
and (n995, n992, n994);
xnor (n995_xnor, n995, n995);
xor (n996, n948_mux, n949_mux);
xor (n996, n948, n949);
xnor (n996_xnor, n996, n996);
and (n997, n994_mux, n996_mux);
and (n997, n994, n996);
xnor (n997_xnor, n997, n997);
and (n998, n992_mux, n996_mux);
and (n998, n992, n996);
xnor (n998_xnor, n998, n998);
or (n999_1, n997_mux, n998_mux);
or (n999, n995_mux, n999_1);
or (n999_1, n997, n998);
or (n999, n995, n999_1);
xnor (n999_xnor, n999, n999);
xor (n1000, n980_mux, n981_mux);
xor (n1000, n980, n981);
xnor (n1000_xnor, n1000, n1000);
xor (n1001, n1000_mux, n985_mux);
xor (n1001, n1000, n985);
xnor (n1001_xnor, n1001, n1001);
and (n1002, n999_mux, n1001_mux);
and (n1002, n999, n1001);
xnor (n1002_xnor, n1002, n1002);
xor (n1003, n947_mux, n950_mux);
xor (n1003, n947, n950);
xnor (n1003_xnor, n1003, n1003);
xor (n1004, n1003_mux, n953_mux);
xor (n1004, n1003, n953);
xnor (n1004_xnor, n1004, n1004);
and (n1005, n1001_mux, n1004_mux);
and (n1005, n1001, n1004);
xnor (n1005_xnor, n1005, n1005);
and (n1006, n999_mux, n1004_mux);
and (n1006, n999, n1004);
xnor (n1006_xnor, n1006, n1006);
or (n1007_1, n1005_mux, n1006_mux);
or (n1007, n1002_mux, n1007_1);
or (n1007_1, n1005, n1006);
or (n1007, n1002, n1007_1);
xnor (n1007_xnor, n1007, n1007);
and (n1008, n988_mux, n1007_mux);
and (n1008, n988, n1007);
xnor (n1008_xnor, n1008, n1008);
xor (n1009, n956_mux, n958_mux);
xor (n1009, n956, n958);
xnor (n1009_xnor, n1009, n1009);
xor (n1010, n1009_mux, n961_mux);
xor (n1010, n1009, n961);
xnor (n1010_xnor, n1010, n1010);
and (n1011, n1007_mux, n1010_mux);
and (n1011, n1007, n1010);
xnor (n1011_xnor, n1011, n1011);
and (n1012, n988_mux, n1010_mux);
and (n1012, n988, n1010);
xnor (n1012_xnor, n1012, n1012);
or (n1013_1, n1011_mux, n1012_mux);
or (n1013, n1008_mux, n1013_1);
or (n1013_1, n1011, n1012);
or (n1013, n1008, n1013_1);
xnor (n1013_xnor, n1013, n1013);
and (n1014, n977_mux, n1013_mux);
and (n1014, n977, n1013);
xnor (n1014_xnor, n1014, n1014);
xor (n1015, n977_mux, n1013_mux);
xor (n1015, n977, n1013);
xnor (n1015_xnor, n1015, n1015);
xor (n1016, n988_mux, n1007_mux);
xor (n1016, n988, n1007);
xnor (n1016_xnor, n1016, n1016);
xor (n1017, n1016_mux, n1010_mux);
xor (n1017, n1016, n1010);
xnor (n1017_xnor, n1017, n1017);
and (n531, n474_mux, n472_mux);
and (n531, n474, n472);
xnor (n531_xnor, n531, n531);
and (n532, n478_mux, n475_mux);
and (n532, n478, n475);
xnor (n532_xnor, n532, n532);
and (n1018, n531_mux, n532_mux);
and (n1018, n531, n532);
xnor (n1018_xnor, n1018, n1018);
and (n534, n486_mux, n479_mux);
and (n534, n486, n479);
xnor (n534_xnor, n534, n534);
and (n1019, n532_mux, n534_mux);
and (n1019, n532, n534);
xnor (n1019_xnor, n1019, n1019);
and (n1020, n531_mux, n534_mux);
and (n1020, n531, n534);
xnor (n1020_xnor, n1020, n1020);
or (n1021_1, n1019_mux, n1020_mux);
or (n1021, n1018_mux, n1021_1);
or (n1021_1, n1019, n1020);
or (n1021, n1018, n1021_1);
xnor (n1021_xnor, n1021, n1021);
not(n1022, n474_mux);
not(n1022, n474);
xnor (n1022_xnor, n1022, n1022);
and (n1023, n546_mux, n474_mux);
and (n1023, n546, n474);
xnor (n1023_xnor, n1023, n1023);
nor (n1024, n1022_mux, n1023_mux);
nor (n1024, n1022, n1023);
xnor (n1024_xnor, n1024, n1024);
and (n1025, n1021_mux, n1024_mux);
and (n1025, n1021, n1024);
xnor (n1025_xnor, n1025, n1025);
and (n1026, n550_mux, n487_mux);
and (n1026, n550, n487);
xnor (n1026_xnor, n1026, n1026);
not(n1027, n487_mux);
not(n1027, n487);
xnor (n1027_xnor, n1027, n1027);
nor (n1028, n1026_mux, n1027_mux);
nor (n1028, n1026, n1027);
xnor (n1028_xnor, n1028, n1028);
and (n1029, n1024_mux, n1028_mux);
and (n1029, n1024, n1028);
xnor (n1029_xnor, n1029, n1029);
and (n1030, n1021_mux, n1028_mux);
and (n1030, n1021, n1028);
xnor (n1030_xnor, n1030, n1030);
or (n1031_1, n1029_mux, n1030_mux);
or (n1031, n1025_mux, n1031_1);
or (n1031_1, n1029, n1030);
or (n1031, n1025, n1031_1);
xnor (n1031_xnor, n1031, n1031);
and (n527, n512_mux, n513_mux);
and (n527, n512, n513);
xnor (n527_xnor, n527, n527);
and (n528, n513_mux, n516_mux);
and (n528, n513, n516);
xnor (n528_xnor, n528, n528);
and (n529, n512_mux, n516_mux);
and (n529, n512, n516);
xnor (n529_xnor, n529, n529);
or (n530_1, n528_mux, n529_mux);
or (n530, n527_mux, n530_1);
or (n530_1, n528, n529);
or (n530, n527, n530_1);
xnor (n530_xnor, n530, n530);
xor (n533, n531_mux, n532_mux);
xor (n533, n531, n532);
xnor (n533_xnor, n533, n533);
xor (n535, n533_mux, n534_mux);
xor (n535, n533, n534);
xnor (n535_xnor, n535, n535);
and (n1032, n530_mux, n535_mux);
and (n1032, n530, n535);
xnor (n1032_xnor, n1032, n1032);
xor (n539, n537_mux, n538_mux);
xor (n539, n537, n538);
xnor (n539_xnor, n539, n539);
xor (n541, n539_mux, n540_mux);
xor (n541, n539, n540);
xnor (n541_xnor, n541, n541);
and (n1033, n535_mux, n541_mux);
and (n1033, n535, n541);
xnor (n1033_xnor, n1033, n1033);
and (n1034, n530_mux, n541_mux);
and (n1034, n530, n541);
xnor (n1034_xnor, n1034, n1034);
or (n1035_1, n1033_mux, n1034_mux);
or (n1035, n1032_mux, n1035_1);
or (n1035_1, n1033, n1034);
or (n1035, n1032, n1035_1);
xnor (n1035_xnor, n1035, n1035);
xor (n1036, n1021_mux, n1024_mux);
xor (n1036, n1021, n1024);
xnor (n1036_xnor, n1036, n1036);
xor (n1037, n1036_mux, n1028_mux);
xor (n1037, n1036, n1028);
xnor (n1037_xnor, n1037, n1037);
and (n1038, n1035_mux, n1037_mux);
and (n1038, n1035, n1037);
xnor (n1038_xnor, n1038, n1038);
xor (n1039, n992_mux, n994_mux);
xor (n1039, n992, n994);
xnor (n1039_xnor, n1039, n1039);
xor (n1040, n1039_mux, n996_mux);
xor (n1040, n1039, n996);
xnor (n1040_xnor, n1040, n1040);
and (n1041, n1037_mux, n1040_mux);
and (n1041, n1037, n1040);
xnor (n1041_xnor, n1041, n1041);
and (n1042, n1035_mux, n1040_mux);
and (n1042, n1035, n1040);
xnor (n1042_xnor, n1042, n1042);
or (n1043_1, n1041_mux, n1042_mux);
or (n1043, n1038_mux, n1043_1);
or (n1043_1, n1041, n1042);
or (n1043, n1038, n1043_1);
xnor (n1043_xnor, n1043, n1043);
and (n1044, n1031_mux, n1043_mux);
and (n1044, n1031, n1043);
xnor (n1044_xnor, n1044, n1044);
xor (n1045, n999_mux, n1001_mux);
xor (n1045, n999, n1001);
xnor (n1045_xnor, n1045, n1045);
xor (n1046, n1045_mux, n1004_mux);
xor (n1046, n1045, n1004);
xnor (n1046_xnor, n1046, n1046);
and (n1047, n1043_mux, n1046_mux);
and (n1047, n1043, n1046);
xnor (n1047_xnor, n1047, n1047);
and (n1048, n1031_mux, n1046_mux);
and (n1048, n1031, n1046);
xnor (n1048_xnor, n1048, n1048);
or (n1049_1, n1047_mux, n1048_mux);
or (n1049, n1044_mux, n1049_1);
or (n1049_1, n1047, n1048);
or (n1049, n1044, n1049_1);
xnor (n1049_xnor, n1049, n1049);
and (n1050, n1017_mux, n1049_mux);
and (n1050, n1017, n1049);
xnor (n1050_xnor, n1050, n1050);
xor (n1051, n1017_mux, n1049_mux);
xor (n1051, n1017, n1049);
xnor (n1051_xnor, n1051, n1051);
xor (n1052, n1031_mux, n1043_mux);
xor (n1052, n1031, n1043);
xnor (n1052_xnor, n1052, n1052);
xor (n1053, n1052_mux, n1046_mux);
xor (n1053, n1052, n1046);
xnor (n1053_xnor, n1053, n1053);
not(n544, n471_mux);
not(n544, n471);
xnor (n544_xnor, n544, n544);
and (n547, n546_mux, n471_mux);
and (n547, n546, n471);
xnor (n547_xnor, n547, n547);
nor (n548, n544_mux, n547_mux);
nor (n548, n544, n547);
xnor (n548_xnor, n548, n548);
and (n551, n550_mux, n491_mux);
and (n551, n550, n491);
xnor (n551_xnor, n551, n551);
not(n552, n491_mux);
not(n552, n491);
xnor (n552_xnor, n552, n552);
nor (n553, n551_mux, n552_mux);
nor (n553, n551, n552);
xnor (n553_xnor, n553, n553);
and (n1054, n548_mux, n553_mux);
and (n1054, n548, n553);
xnor (n1054_xnor, n1054, n1054);
and (n523, n508_mux, n510_mux);
and (n523, n508, n510);
xnor (n523_xnor, n523, n523);
and (n524, n510_mux, n517_mux);
and (n524, n510, n517);
xnor (n524_xnor, n524, n524);
and (n525, n508_mux, n517_mux);
and (n525, n508, n517);
xnor (n525_xnor, n525, n525);
or (n526_1, n524_mux, n525_mux);
or (n526, n523_mux, n526_1);
or (n526_1, n524, n525);
or (n526, n523, n526_1);
xnor (n526_xnor, n526, n526);
xor (n536, n530_mux, n535_mux);
xor (n536, n530, n535);
xnor (n536_xnor, n536, n536);
xor (n542, n536_mux, n541_mux);
xor (n542, n536, n541);
xnor (n542_xnor, n542, n542);
and (n1055, n526_mux, n542_mux);
and (n1055, n526, n542);
xnor (n1055_xnor, n1055, n1055);
xor (n554, n548_mux, n553_mux);
xor (n554, n548, n553);
xnor (n554_xnor, n554, n554);
and (n1056, n542_mux, n554_mux);
and (n1056, n542, n554);
xnor (n1056_xnor, n1056, n1056);
and (n1057, n526_mux, n554_mux);
and (n1057, n526, n554);
xnor (n1057_xnor, n1057, n1057);
or (n1058_1, n1056_mux, n1057_mux);
or (n1058, n1055_mux, n1058_1);
or (n1058_1, n1056, n1057);
or (n1058, n1055, n1058_1);
xnor (n1058_xnor, n1058, n1058);
and (n1059, n1054_mux, n1058_mux);
and (n1059, n1054, n1058);
xnor (n1059_xnor, n1059, n1059);
xor (n1060, n1035_mux, n1037_mux);
xor (n1060, n1035, n1037);
xnor (n1060_xnor, n1060, n1060);
xor (n1061, n1060_mux, n1040_mux);
xor (n1061, n1060, n1040);
xnor (n1061_xnor, n1061, n1061);
and (n1062, n1058_mux, n1061_mux);
and (n1062, n1058, n1061);
xnor (n1062_xnor, n1062, n1062);
and (n1063, n1054_mux, n1061_mux);
and (n1063, n1054, n1061);
xnor (n1063_xnor, n1063, n1063);
or (n1064_1, n1062_mux, n1063_mux);
or (n1064, n1059_mux, n1064_1);
or (n1064_1, n1062, n1063);
or (n1064, n1059, n1064_1);
xnor (n1064_xnor, n1064, n1064);
and (n1065, n1053_mux, n1064_mux);
and (n1065, n1053, n1064);
xnor (n1065_xnor, n1065, n1065);
xor (n1066, n1053_mux, n1064_mux);
xor (n1066, n1053, n1064);
xnor (n1066_xnor, n1066, n1066);
xor (n1067, n1054_mux, n1058_mux);
xor (n1067, n1054, n1058);
xnor (n1067_xnor, n1067, n1067);
xor (n1068, n1067_mux, n1061_mux);
xor (n1068, n1067, n1061);
xnor (n1068_xnor, n1068, n1068);
and (n477, n473_mux, n476_mux);
and (n477, n473, n476);
xnor (n477_xnor, n477, n477);
and (n481, n476_mux, n480_mux);
and (n481, n476, n480);
xnor (n481_xnor, n481, n481);
and (n482, n473_mux, n480_mux);
and (n482, n473, n480);
xnor (n482_xnor, n482, n482);
or (n483_1, n481_mux, n482_mux);
or (n483, n477_mux, n483_1);
or (n483_1, n481, n482);
or (n483, n477, n483_1);
xnor (n483_xnor, n483, n483);
and (n507, n504_mux, n506_mux);
and (n507, n504, n506);
xnor (n507_xnor, n507, n507);
and (n519, n506_mux, n518_mux);
and (n519, n506, n518);
xnor (n519_xnor, n519, n519);
and (n520, n504_mux, n518_mux);
and (n520, n504, n518);
xnor (n520_xnor, n520, n520);
or (n521_1, n519_mux, n520_mux);
or (n521, n507_mux, n521_1);
or (n521_1, n519, n520);
or (n521, n507, n521_1);
xnor (n521_xnor, n521, n521);
and (n1069, n483_mux, n521_mux);
and (n1069, n483, n521);
xnor (n1069_xnor, n1069, n1069);
xor (n543, n526_mux, n542_mux);
xor (n543, n526, n542);
xnor (n543_xnor, n543, n543);
xor (n555, n543_mux, n554_mux);
xor (n555, n543, n554);
xnor (n555_xnor, n555, n555);
and (n1070, n521_mux, n555_mux);
and (n1070, n521, n555);
xnor (n1070_xnor, n1070, n1070);
and (n1071, n483_mux, n555_mux);
and (n1071, n483, n555);
xnor (n1071_xnor, n1071, n1071);
or (n1072_1, n1070_mux, n1071_mux);
or (n1072, n1069_mux, n1072_1);
or (n1072_1, n1070, n1071);
or (n1072, n1069, n1072_1);
xnor (n1072_xnor, n1072, n1072);
and (n1073, n1068_mux, n1072_mux);
and (n1073, n1068, n1072);
xnor (n1073_xnor, n1073, n1073);
xor (n1074, n1068_mux, n1072_mux);
xor (n1074, n1068, n1072);
xnor (n1074_xnor, n1074, n1074);
xor (n522, n483_mux, n521_mux);
xor (n522, n483, n521);
xnor (n522_xnor, n522, n522);
xor (n556, n522_mux, n555_mux);
xor (n556, n522, n555);
xnor (n556_xnor, n556, n556);
and (n581, n559_mux, n580_mux);
and (n581, n559, n580);
xnor (n581_xnor, n581, n581);
and (n584, n580_mux, n583_mux);
and (n584, n580, n583);
xnor (n584_xnor, n584, n584);
and (n585, n559_mux, n583_mux);
and (n585, n559, n583);
xnor (n585_xnor, n585, n585);
or (n586_1, n584_mux, n585_mux);
or (n586, n581_mux, n586_1);
or (n586_1, n584, n585);
or (n586, n581, n586_1);
xnor (n586_xnor, n586, n586);
and (n1075, n556_mux, n586_mux);
and (n1075, n556, n586);
xnor (n1075_xnor, n1075, n1075);
xor (n587, n556_mux, n586_mux);
xor (n587, n556, n586);
xnor (n587_xnor, n587, n587);
and (n614, n589_mux, n613_mux);
and (n614, n589, n613);
xnor (n614_xnor, n614, n614);
and (n634, n615_mux, n633_mux);
and (n634, n615, n633);
xnor (n634_xnor, n634, n634);
or (n635, n614_mux, n634_mux);
or (n635, n614, n634);
xnor (n635_xnor, n635, n635);
and (n1076, n587_mux, n635_mux);
and (n1076, n587, n635);
xnor (n1076_xnor, n1076, n1076);
or (n1077, n1075_mux, n1076_mux);
or (n1077, n1075, n1076);
xnor (n1077_xnor, n1077, n1077);
and (n1078, n1074_mux, n1077_mux);
and (n1078, n1074, n1077);
xnor (n1078_xnor, n1078, n1078);
or (n1079, n1073_mux, n1078_mux);
or (n1079, n1073, n1078);
xnor (n1079_xnor, n1079, n1079);
and (n1080, n1066_mux, n1079_mux);
and (n1080, n1066, n1079);
xnor (n1080_xnor, n1080, n1080);
or (n1081, n1065_mux, n1080_mux);
or (n1081, n1065, n1080);
xnor (n1081_xnor, n1081, n1081);
and (n1082, n1051_mux, n1081_mux);
and (n1082, n1051, n1081);
xnor (n1082_xnor, n1082, n1082);
or (n1083, n1050_mux, n1082_mux);
or (n1083, n1050, n1082);
xnor (n1083_xnor, n1083, n1083);
and (n1084, n1015_mux, n1083_mux);
and (n1084, n1015, n1083);
xnor (n1084_xnor, n1084, n1084);
or (n1085, n1014_mux, n1084_mux);
or (n1085, n1014, n1084);
xnor (n1085_xnor, n1085, n1085);
and (n1086, n975_mux, n1085_mux);
and (n1086, n975, n1085);
xnor (n1086_xnor, n1086, n1086);
or (n1087, n974_mux, n1086_mux);
or (n1087, n974, n1086);
xnor (n1087_xnor, n1087, n1087);
and (n1088, n938_mux, n1087_mux);
and (n1088, n938, n1087);
xnor (n1088_xnor, n1088, n1088);
or (n1089, n937_mux, n1088_mux);
or (n1089, n937, n1088);
xnor (n1089_xnor, n1089, n1089);
and (n1090, n895_mux, n1089_mux);
and (n1090, n895, n1089);
xnor (n1090_xnor, n1090, n1090);
or (n1091, n894_mux, n1090_mux);
or (n1091, n894, n1090);
xnor (n1091_xnor, n1091, n1091);
buf(n1092, n1091_mux);
buf(n1092, n1091);
xnor (n1092_xnor, n1092, n1092);
buf(n1357, n1092_mux);
buf(n1357, n1092);
xnor (n1357_xnor, n1357, n1357);
xor (n1093, n895_mux, n1089_mux);
xor (n1093, n895, n1089);
xnor (n1093_xnor, n1093, n1093);
buf(n1094, n1093_mux);
buf(n1094, n1093);
xnor (n1094_xnor, n1094, n1094);
buf(n1358, n1094_mux);
buf(n1358, n1094);
xnor (n1358_xnor, n1358, n1358);
xor (n1095, n938_mux, n1087_mux);
xor (n1095, n938, n1087);
xnor (n1095_xnor, n1095, n1095);
buf(n1096, n1095_mux);
buf(n1096, n1095);
xnor (n1096_xnor, n1096, n1096);
buf(n1359, n1096_mux);
buf(n1359, n1096);
xnor (n1359_xnor, n1359, n1359);
xor (n1097, n975_mux, n1085_mux);
xor (n1097, n975, n1085);
xnor (n1097_xnor, n1097, n1097);
buf(n1098, n1097_mux);
buf(n1098, n1097);
xnor (n1098_xnor, n1098, n1098);
buf(n1360, n1098_mux);
buf(n1360, n1098);
xnor (n1360_xnor, n1360, n1360);
xor (n1099, n1015_mux, n1083_mux);
xor (n1099, n1015, n1083);
xnor (n1099_xnor, n1099, n1099);
buf(n1100, n1099_mux);
buf(n1100, n1099);
xnor (n1100_xnor, n1100, n1100);
buf(n1361, n1100_mux);
buf(n1361, n1100);
xnor (n1361_xnor, n1361, n1361);
xor (n1101, n1051_mux, n1081_mux);
xor (n1101, n1051, n1081);
xnor (n1101_xnor, n1101, n1101);
buf(n1102, n1101_mux);
buf(n1102, n1101);
xnor (n1102_xnor, n1102, n1102);
buf(n1362, n1102_mux);
buf(n1362, n1102);
xnor (n1362_xnor, n1362, n1362);
xor (n1103, n1066_mux, n1079_mux);
xor (n1103, n1066, n1079);
xnor (n1103_xnor, n1103, n1103);
buf(n1104, n1103_mux);
buf(n1104, n1103);
xnor (n1104_xnor, n1104, n1104);
buf(n1363, n1104_mux);
buf(n1363, n1104);
xnor (n1363_xnor, n1363, n1363);
buf(n1348, n845_mux);
buf(n1348, n845);
xnor (n1348_xnor, n1348, n1348);
xor (n1105, n1074_mux, n1077_mux);
xor (n1105, n1074, n1077);
xnor (n1105_xnor, n1105, n1105);
buf(n1106, n1105_mux);
buf(n1106, n1105);
xnor (n1106_xnor, n1106, n1106);
buf(n1364, n1106_mux);
buf(n1364, n1106);
xnor (n1364_xnor, n1364, n1364);
and (n1373, n1348_mux, n1364_mux);
and (n1373, n1348, n1364);
xnor (n1373_xnor, n1373, n1373);
buf(n1349, n834_mux);
buf(n1349, n834);
xnor (n1349_xnor, n1349, n1349);
xor (n636, n587_mux, n635_mux);
xor (n636, n587, n635);
xnor (n636_xnor, n636, n636);
buf(n637, n636_mux);
buf(n637, n636);
xnor (n637_xnor, n637, n637);
buf(n1365, n637_mux);
buf(n1365, n637);
xnor (n1365_xnor, n1365, n1365);
and (n1374, n1349_mux, n1365_mux);
and (n1374, n1349, n1365);
xnor (n1374_xnor, n1374, n1374);
buf(n1350, n815_mux);
buf(n1350, n815);
xnor (n1350_xnor, n1350, n1350);
buf(n1366, n642_mux);
buf(n1366, n642);
xnor (n1366_xnor, n1366, n1366);
and (n1375, n1350_mux, n1366_mux);
and (n1375, n1350, n1366);
xnor (n1375_xnor, n1375, n1375);
buf(n1351, n796_mux);
buf(n1351, n796);
xnor (n1351_xnor, n1351, n1351);
buf(n1367, n649_mux);
buf(n1367, n649);
xnor (n1367_xnor, n1367, n1367);
and (n1376, n1351_mux, n1367_mux);
and (n1376, n1351, n1367);
xnor (n1376_xnor, n1376, n1376);
buf(n1352, n777_mux);
buf(n1352, n777);
xnor (n1352_xnor, n1352, n1352);
buf(n1368, n656_mux);
buf(n1368, n656);
xnor (n1368_xnor, n1368, n1368);
and (n1377, n1352_mux, n1368_mux);
and (n1377, n1352, n1368);
xnor (n1377_xnor, n1377, n1377);
buf(n1353, n758_mux);
buf(n1353, n758);
xnor (n1353_xnor, n1353, n1353);
buf(n1369, n663_mux);
buf(n1369, n663);
xnor (n1369_xnor, n1369, n1369);
and (n1378, n1353_mux, n1369_mux);
and (n1378, n1353, n1369);
xnor (n1378_xnor, n1378, n1378);
buf(n1354, n739_mux);
buf(n1354, n739);
xnor (n1354_xnor, n1354, n1354);
buf(n1370, n670_mux);
buf(n1370, n670);
xnor (n1370_xnor, n1370, n1370);
and (n1379, n1354_mux, n1370_mux);
and (n1379, n1354, n1370);
xnor (n1379_xnor, n1379, n1379);
buf(n1355, n720_mux);
buf(n1355, n720);
xnor (n1355_xnor, n1355, n1355);
buf(n1371, n677_mux);
buf(n1371, n677);
xnor (n1371_xnor, n1371, n1371);
and (n1380, n1355_mux, n1371_mux);
and (n1380, n1355, n1371);
xnor (n1380_xnor, n1380, n1380);
buf(n1356, n707_mux);
buf(n1356, n707);
xnor (n1356_xnor, n1356, n1356);
buf(n1372, n684_mux);
buf(n1372, n684);
xnor (n1372_xnor, n1372, n1372);
and (n1381, n1356_mux, n1372_mux);
and (n1381, n1356, n1372);
xnor (n1381_xnor, n1381, n1381);
and (n1382, n1371_mux, n1381_mux);
and (n1382, n1371, n1381);
xnor (n1382_xnor, n1382, n1382);
and (n1383, n1355_mux, n1381_mux);
and (n1383, n1355, n1381);
xnor (n1383_xnor, n1383, n1383);
or (n1384_1, n1382_mux, n1383_mux);
or (n1384, n1380_mux, n1384_1);
or (n1384_1, n1382, n1383);
or (n1384, n1380, n1384_1);
xnor (n1384_xnor, n1384, n1384);
and (n1385, n1370_mux, n1384_mux);
and (n1385, n1370, n1384);
xnor (n1385_xnor, n1385, n1385);
and (n1386, n1354_mux, n1384_mux);
and (n1386, n1354, n1384);
xnor (n1386_xnor, n1386, n1386);
or (n1387_1, n1385_mux, n1386_mux);
or (n1387, n1379_mux, n1387_1);
or (n1387_1, n1385, n1386);
or (n1387, n1379, n1387_1);
xnor (n1387_xnor, n1387, n1387);
and (n1388, n1369_mux, n1387_mux);
and (n1388, n1369, n1387);
xnor (n1388_xnor, n1388, n1388);
and (n1389, n1353_mux, n1387_mux);
and (n1389, n1353, n1387);
xnor (n1389_xnor, n1389, n1389);
or (n1390_1, n1388_mux, n1389_mux);
or (n1390, n1378_mux, n1390_1);
or (n1390_1, n1388, n1389);
or (n1390, n1378, n1390_1);
xnor (n1390_xnor, n1390, n1390);
and (n1391, n1368_mux, n1390_mux);
and (n1391, n1368, n1390);
xnor (n1391_xnor, n1391, n1391);
and (n1392, n1352_mux, n1390_mux);
and (n1392, n1352, n1390);
xnor (n1392_xnor, n1392, n1392);
or (n1393_1, n1391_mux, n1392_mux);
or (n1393, n1377_mux, n1393_1);
or (n1393_1, n1391, n1392);
or (n1393, n1377, n1393_1);
xnor (n1393_xnor, n1393, n1393);
and (n1394, n1367_mux, n1393_mux);
and (n1394, n1367, n1393);
xnor (n1394_xnor, n1394, n1394);
and (n1395, n1351_mux, n1393_mux);
and (n1395, n1351, n1393);
xnor (n1395_xnor, n1395, n1395);
or (n1396_1, n1394_mux, n1395_mux);
or (n1396, n1376_mux, n1396_1);
or (n1396_1, n1394, n1395);
or (n1396, n1376, n1396_1);
xnor (n1396_xnor, n1396, n1396);
and (n1397, n1366_mux, n1396_mux);
and (n1397, n1366, n1396);
xnor (n1397_xnor, n1397, n1397);
and (n1398, n1350_mux, n1396_mux);
and (n1398, n1350, n1396);
xnor (n1398_xnor, n1398, n1398);
or (n1399_1, n1397_mux, n1398_mux);
or (n1399, n1375_mux, n1399_1);
or (n1399_1, n1397, n1398);
or (n1399, n1375, n1399_1);
xnor (n1399_xnor, n1399, n1399);
and (n1400, n1365_mux, n1399_mux);
and (n1400, n1365, n1399);
xnor (n1400_xnor, n1400, n1400);
and (n1401, n1349_mux, n1399_mux);
and (n1401, n1349, n1399);
xnor (n1401_xnor, n1401, n1401);
or (n1402_1, n1400_mux, n1401_mux);
or (n1402, n1374_mux, n1402_1);
or (n1402_1, n1400, n1401);
or (n1402, n1374, n1402_1);
xnor (n1402_xnor, n1402, n1402);
and (n1403, n1364_mux, n1402_mux);
and (n1403, n1364, n1402);
xnor (n1403_xnor, n1403, n1403);
and (n1404, n1348_mux, n1402_mux);
and (n1404, n1348, n1402);
xnor (n1404_xnor, n1404, n1404);
or (n1405_1, n1403_mux, n1404_mux);
or (n1405, n1373_mux, n1405_1);
or (n1405_1, n1403, n1404);
or (n1405, n1373, n1405_1);
xnor (n1405_xnor, n1405, n1405);
and (n1406, n1363_mux, n1405_mux);
and (n1406, n1363, n1405);
xnor (n1406_xnor, n1406, n1406);
and (n1407, n1362_mux, n1406_mux);
and (n1407, n1362, n1406);
xnor (n1407_xnor, n1407, n1407);
and (n1408, n1361_mux, n1407_mux);
and (n1408, n1361, n1407);
xnor (n1408_xnor, n1408, n1408);
and (n1409, n1360_mux, n1408_mux);
and (n1409, n1360, n1408);
xnor (n1409_xnor, n1409, n1409);
and (n1410, n1359_mux, n1409_mux);
and (n1410, n1359, n1409);
xnor (n1410_xnor, n1410, n1410);
and (n1411, n1358_mux, n1410_mux);
and (n1411, n1358, n1410);
xnor (n1411_xnor, n1411, n1411);
and (n1412, n1357_mux, n1411_mux);
and (n1412, n1357, n1411);
xnor (n1412_xnor, n1412, n1412);
buf(n1413, n1412_mux);
buf(n1413, n1412);
xnor (n1413_xnor, n1413, n1413);
buf(n163, n1413_mux);
buf(g144, n163);
buf(n163, n1413);
buf(g144, n163);
xnor (g144_xnor, g144, g144);
xor (n1414, n1357_mux, n1411_mux);
xor (n1414, n1357, n1411);
xnor (n1414_xnor, n1414, n1414);
buf(n1415, n1414_mux);
buf(n1415, n1414);
xnor (n1415_xnor, n1415, n1415);
buf(n164, n1415_mux);
buf(g145, n164);
buf(n164, n1415);
buf(g145, n164);
xnor (g145_xnor, g145, g145);
xor (n1416, n1358_mux, n1410_mux);
xor (n1416, n1358, n1410);
xnor (n1416_xnor, n1416, n1416);
buf(n1417, n1416_mux);
buf(n1417, n1416);
xnor (n1417_xnor, n1417, n1417);
buf(n165, n1417_mux);
buf(g146, n165);
buf(n165, n1417);
buf(g146, n165);
xnor (g146_xnor, g146, g146);
xor (n1418, n1359_mux, n1409_mux);
xor (n1418, n1359, n1409);
xnor (n1418_xnor, n1418, n1418);
buf(n1419, n1418_mux);
buf(n1419, n1418);
xnor (n1419_xnor, n1419, n1419);
buf(n166, n1419_mux);
buf(g147, n166);
buf(n166, n1419);
buf(g147, n166);
xnor (g147_xnor, g147, g147);
xor (n1420, n1360_mux, n1408_mux);
xor (n1420, n1360, n1408);
xnor (n1420_xnor, n1420, n1420);
buf(n1421, n1420_mux);
buf(n1421, n1420);
xnor (n1421_xnor, n1421, n1421);
buf(n167, n1421_mux);
buf(g148, n167);
buf(n167, n1421);
buf(g148, n167);
xnor (g148_xnor, g148, g148);
xor (n1422, n1361_mux, n1407_mux);
xor (n1422, n1361, n1407);
xnor (n1422_xnor, n1422, n1422);
buf(n1423, n1422_mux);
buf(n1423, n1422);
xnor (n1423_xnor, n1423, n1423);
buf(n168, n1423_mux);
buf(g149, n168);
buf(n168, n1423);
buf(g149, n168);
xnor (g149_xnor, g149, g149);
xor (n1424, n1362_mux, n1406_mux);
xor (n1424, n1362, n1406);
xnor (n1424_xnor, n1424, n1424);
buf(n1425, n1424_mux);
buf(n1425, n1424);
xnor (n1425_xnor, n1425, n1425);
buf(n169, n1425_mux);
buf(g150, n169);
buf(n169, n1425);
buf(g150, n169);
xnor (g150_xnor, g150, g150);
xor (n1426, n1363_mux, n1405_mux);
xor (n1426, n1363, n1405);
xnor (n1426_xnor, n1426, n1426);
buf(n1427, n1426_mux);
buf(n1427, n1426);
xnor (n1427_xnor, n1427, n1427);
buf(n170, n1427_mux);
buf(g151, n170);
buf(n170, n1427);
buf(g151, n170);
xnor (g151_xnor, g151, g151);
xor (n1428, n1348_mux, n1364_mux);
xor (n1428, n1348, n1364);
xnor (n1428_xnor, n1428, n1428);
xor (n1429, n1428_mux, n1402_mux);
xor (n1429, n1428, n1402);
xnor (n1429_xnor, n1429, n1429);
buf(n1430, n1429_mux);
buf(n1430, n1429);
xnor (n1430_xnor, n1430, n1430);
buf(n171, n1430_mux);
buf(g152, n171);
buf(n171, n1430);
buf(g152, n171);
xnor (g152_xnor, g152, g152);
xor (n1431, n1349_mux, n1365_mux);
xor (n1431, n1349, n1365);
xnor (n1431_xnor, n1431, n1431);
xor (n1432, n1431_mux, n1399_mux);
xor (n1432, n1431, n1399);
xnor (n1432_xnor, n1432, n1432);
buf(n1433, n1432_mux);
buf(n1433, n1432);
xnor (n1433_xnor, n1433, n1433);
buf(n172, n1433_mux);
buf(g153, n172);
buf(n172, n1433);
buf(g153, n172);
xnor (g153_xnor, g153, g153);
xor (n1434, n1350_mux, n1366_mux);
xor (n1434, n1350, n1366);
xnor (n1434_xnor, n1434, n1434);
xor (n1435, n1434_mux, n1396_mux);
xor (n1435, n1434, n1396);
xnor (n1435_xnor, n1435, n1435);
buf(n1436, n1435_mux);
buf(n1436, n1435);
xnor (n1436_xnor, n1436, n1436);
buf(n173, n1436_mux);
buf(g154, n173);
buf(n173, n1436);
buf(g154, n173);
xnor (g154_xnor, g154, g154);
xor (n1437, n1351_mux, n1367_mux);
xor (n1437, n1351, n1367);
xnor (n1437_xnor, n1437, n1437);
xor (n1438, n1437_mux, n1393_mux);
xor (n1438, n1437, n1393);
xnor (n1438_xnor, n1438, n1438);
buf(n1439, n1438_mux);
buf(n1439, n1438);
xnor (n1439_xnor, n1439, n1439);
buf(n174, n1439_mux);
buf(g155, n174);
buf(n174, n1439);
buf(g155, n174);
xnor (g155_xnor, g155, g155);
xor (n1440, n1352_mux, n1368_mux);
xor (n1440, n1352, n1368);
xnor (n1440_xnor, n1440, n1440);
xor (n1441, n1440_mux, n1390_mux);
xor (n1441, n1440, n1390);
xnor (n1441_xnor, n1441, n1441);
buf(n1442, n1441_mux);
buf(n1442, n1441);
xnor (n1442_xnor, n1442, n1442);
buf(n175, n1442_mux);
buf(g156, n175);
buf(n175, n1442);
buf(g156, n175);
xnor (g156_xnor, g156, g156);
xor (n1443, n1353_mux, n1369_mux);
xor (n1443, n1353, n1369);
xnor (n1443_xnor, n1443, n1443);
xor (n1444, n1443_mux, n1387_mux);
xor (n1444, n1443, n1387);
xnor (n1444_xnor, n1444, n1444);
buf(n1445, n1444_mux);
buf(n1445, n1444);
xnor (n1445_xnor, n1445, n1445);
buf(n176, n1445_mux);
buf(g157, n176);
buf(n176, n1445);
buf(g157, n176);
xnor (g157_xnor, g157, g157);
xor (n1446, n1354_mux, n1370_mux);
xor (n1446, n1354, n1370);
xnor (n1446_xnor, n1446, n1446);
xor (n1447, n1446_mux, n1384_mux);
xor (n1447, n1446, n1384);
xnor (n1447_xnor, n1447, n1447);
buf(n1448, n1447_mux);
buf(n1448, n1447);
xnor (n1448_xnor, n1448, n1448);
buf(n177, n1448_mux);
buf(g158, n177);
buf(n177, n1448);
buf(g158, n177);
xnor (g158_xnor, g158, g158);
xor (n1449, n1355_mux, n1371_mux);
xor (n1449, n1355, n1371);
xnor (n1449_xnor, n1449, n1449);
xor (n1450, n1449_mux, n1381_mux);
xor (n1450, n1449, n1381);
xnor (n1450_xnor, n1450, n1450);
buf(n1451, n1450_mux);
buf(n1451, n1450);
xnor (n1451_xnor, n1451, n1451);
buf(n178, n1451_mux);
buf(g159, n178);
buf(n178, n1451);
buf(g159, n178);
xnor (g159_xnor, g159, g159);
xor (n1452, n1356_mux, n1372_mux);
xor (n1452, n1356, n1372);
xnor (n1452_xnor, n1452, n1452);
buf(n1453, n1452_mux);
buf(n1453, n1452);
xnor (n1453_xnor, n1453, n1453);
buf(n179, n1453_mux);
buf(g160, n179);
buf(n179, n1453);
buf(g160, n179);
xnor (g160_xnor, g160, g160);
patch p0 (.1'b0(t_0), 
endmodule