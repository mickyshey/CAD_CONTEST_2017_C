module patch (w684, g0, g1, g2, g3, g4, g5, g6, g7);g8, g9, g10, 
input g0, g1, g2, g3, g4, g5, g6, g7;g8, g9, g10, 
output w684;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684;
or (w0, g1, g5);
and (w1, g1, g1);
and (w2, g1, g1);
and (w3, g8, g9);
and (w4, g9, g8);
or (w5, w4, w3);
and (w6, w5, g1);
or (w7, w6, w2);
or (w8, w7, w1);
or (w9, w8, g5);
or (w10, w9, g5);
and (w11, w10, w0);
or (w12, w11, g6);
or (w13, w12, g6);
and (w14, g2, g2);
or (w15, w14, g1);
and (w16, w15, g1);
and (w17, g2, g2);
or (w18, w17, g1);
and (w19, w18, g1);
or (w20, g2, g5);
and (w21, w20, g2);
and (w22, w21, g5);
or (w23, w22, g1);
and (w24, w23, g1);
and (w25, g2, g2);
or (w26, w25, g5);
and (w27, w26, g5);
or (w28, w27, g1);
and (w29, w28, g1);
and (w30, g2, g5);
and (w31, w30, g1);
or (w32, w31, g6);
or (w33, w29, w32);
or (w34, w33, w24);
or (w35, w34, g6);
or (w36, w35, g6);
and (w37, g2, g2);
or (w38, g5, g2);
and (w39, w38, g5);
and (w40, w39, g2);
or (w41, w40, g1);
and (w42, w41, g1);
and (w43, w0, g2);
and (w44, w43, g5);
or (w45, g8, g9);
or (w46, g8, g9);
and (w47, w46, w45);
or (w48, g7, g3);
and (w49, w48, g7);
and (w50, w49, g3);
or (w51, g7, g3);
and (w52, g3, g3);
or (w53, w52, g7);
and (w54, w53, g7);
and (w55, g3, g3);
or (w56, w55, w54);
or (w57, w56, g7);
and (w58, w57, g7);
and (w59, g3, g3);
or (w60, w59, g7);
and (w61, w60, g7);
or (w62, w61, w58);
or (w63, w62, w50);
and (w64, g9, g9);
or (w65, w64, g8);
or (w66, w65, g8);
and (w67, g9, g9);
or (w68, w67, g8);
or (w69, w68, g8);
and (w70, w69, w66);
or (w71, w63, g2);
or (w72, w71, g2);
or (w73, w72, g7);
or (w74, w73, g3);
and (w75, w74, g7);
and (w76, w75, g3);
or (w77, w76, w70);
or (w78, w77, g6);
and (w79, w78, g6);
or (w80, w63, g2);
and (w81, w80, g2);
or (w82, w81, w70);
or (w83, w82, g6);
and (w84, w83, g6);
and (w85, g3, g3);
or (w86, w85, w54);
or (w87, w86, g7);
and (w88, w87, g7);
or (w89, w88, w70);
and (w90, g7, g7);
or (w91, w90, w89);
or (w92, w91, g2);
and (w93, w92, g2);
or (w94, w93, w84);
or (w95, w94, w79);
or (w96, w95, w70);
or (w97, w96, g6);
and (w98, w97, g6);
or (w99, w0, g2);
or (w100, w99, g2);
or (w101, w100, g6);
and (w102, w101, g6);
and (w103, g7, g3);
or (w104, g7, g3);
and (w105, w104, g7);
and (w106, w105, g3);
or (w107, w106, w13);
or (w108, w107, w103);
and (w109, w108, w102);
or (w110, w109, w98);
or (w111, w110, w70);
or (w112, w111, w47);
or (w113, w112, g5);
and (w114, w113, g5);
and (w115, w114, g6);
or (w116, w115, g1);
and (w117, w116, g1);
or (w118, g7, g3);
and (w119, w118, g7);
and (w120, w119, g3);
or (w121, w120, g2);
and (w122, w121, g2);
or (w123, w122, w84);
or (w124, w123, w70);
or (w125, w124, g6);
and (w126, w125, g6);
and (w127, g2, g7);
and (w128, w127, g3);
or (w129, g8, g9);
or (w130, g8, g9);
and (w131, w130, w129);
and (w132, g5, g5);
or (w133, w132, w117);
or (w134, w133, w84);
or (w135, w134, g2);
or (w136, w135, g2);
or (w137, w136, g6);
and (w138, w137, g6);
or (w139, w138, w70);
or (w140, w139, w131);
and (w141, g5, g5);
or (w142, w141, w70);
and (w143, g5, g5);
or (w144, w143, w142);
or (w145, w144, w70);
and (w146, g2, w140);
or (w147, w146, w84);
or (w148, w147, g6);
and (w149, w148, g6);
or (w150, w149, w145);
or (w151, w150, w70);
or (w152, w151, w131);
or (w153, w2, g1);
or (w154, w153, g5);
or (w155, w154, g5);
and (w156, w155, w102);
and (w157, w156, w128);
or (w158, w157, g2);
or (w159, w158, g2);
or (w160, w159, w152);
or (w161, w160, g7);
or (w162, w161, g3);
and (w163, w162, g7);
and (w164, w163, g3);
or (w165, w164, g6);
and (w166, w165, g6);
or (w167, w166, w145);
or (w168, w167, w70);
or (w169, w168, w131);
and (w170, g1, g1);
or (w171, w170, g5);
or (w172, w171, w117);
and (w173, w172, g5);
or (w174, w173, w70);
or (w175, w174, w131);
or (w176, w1, w117);
or (w177, w176, g1);
or (w178, w177, g1);
or (w179, w178, g5);
and (w180, w179, g5);
or (w181, w180, w175);
or (w182, w181, g2);
and (w183, w182, w169);
or (w184, w183, w152);
or (w185, w184, g7);
or (w186, w185, g3);
and (w187, w186, g7);
and (w188, w187, g3);
and (w189, w188, w103);
or (w190, w189, w145);
or (w191, w190, w70);
or (w192, w191, w131);
or (w193, w126, g1);
and (w194, w193, g1);
or (w195, w194, g5);
or (w196, w195, w117);
and (w197, w196, g5);
or (w198, w197, w145);
or (w199, w198, w131);
or (w200, w126, g1);
or (w201, w200, w117);
and (w202, w201, g1);
or (w203, w202, g5);
and (w204, w203, g5);
or (w205, w204, w199);
or (w206, w205, w145);
or (w207, w206, w131);
or (w208, w98, g1);
and (w209, w208, g1);
or (w210, w209, w207);
or (w211, w210, g5);
and (w212, w211, g5);
or (w213, w212, w199);
or (w214, w213, w145);
or (w215, w214, w70);
or (w216, w215, w131);
or (w217, g7, g3);
and (w218, w217, g7);
and (w219, w218, g3);
or (w220, w219, w13);
or (w221, w220, w216);
and (w222, w221, w51);
or (w223, w222, w192);
and (w224, w223, g6);
or (w225, w224, w145);
or (w226, w225, w131);
and (w227, g7, g7);
or (w228, w227, w89);
or (w229, w228, g2);
or (w230, w229, g2);
or (w231, w230, w103);
or (w232, w231, g1);
and (w233, w232, g1);
or (w234, w233, g5);
and (w235, w234, g5);
or (w236, w235, g6);
and (w237, w236, g6);
or (w238, w237, w145);
or (w239, w238, w70);
or (w240, g2, g6);
and (w241, w240, g6);
or (w242, w50, g2);
or (w243, w242, g2);
and (w244, w243, w241);
or (w245, w244, g7);
or (w246, w245, g3);
and (w247, w246, g7);
and (w248, w247, g3);
or (w249, w248, g6);
and (w250, w249, g6);
or (w251, w250, w145);
or (w252, w251, w70);
or (w253, g1, w239);
and (w254, w253, g5);
or (w255, w254, w131);
and (w256, g3, g3);
or (w257, w256, g7);
and (w258, w257, g7);
or (w259, w258, w58);
or (w260, w259, g2);
or (w261, w260, g2);
or (w262, w261, w252);
or (w263, w262, g6);
and (w264, w263, g6);
or (w265, w264, w145);
or (w266, w265, w70);
and (w267, g7, g7);
or (w268, w267, w89);
or (w269, w268, w2);
or (w270, w269, g1);
and (w271, w270, g1);
or (w272, w271, g5);
or (w273, w272, w32);
and (w274, w273, g5);
or (w275, w274, w255);
or (w276, w275, g2);
or (w277, w276, g2);
and (w278, w277, w266);
and (w279, w278, w51);
or (w280, w279, w252);
or (w281, w280, g6);
and (w282, w281, g6);
or (w283, w282, w145);
or (w284, w283, w70);
or (w285, w284, w131);
or (w286, g1, g5);
and (w287, w286, g5);
or (w288, w1, g1);
or (w289, w288, g1);
or (w290, w289, g5);
and (w291, w290, g5);
or (w292, w291, w287);
and (w293, w292, g7);
and (w294, w293, g3);
and (w295, w294, w103);
or (w296, w295, w145);
or (w297, w296, w70);
or (w298, w297, w131);
or (w299, g7, g3);
and (w300, w299, g7);
and (w301, w300, g3);
or (w302, w44, w42);
or (w303, w302, w36);
or (w304, w303, w301);
and (w305, w304, w51);
or (w306, w305, w298);
or (w307, w306, g2);
or (w308, w307, g2);
or (w309, w308, w285);
or (w310, w309, g6);
and (w311, w310, g6);
or (w312, w311, w70);
or (w313, w312, w131);
or (w314, w1, g1);
or (w315, w314, g1);
or (w316, w315, g5);
and (w317, w316, g5);
or (w318, w317, w287);
or (w319, g9, g8);
and (w320, w319, w66);
or (w321, w320, w3);
and (w322, w321, w318);
or (w323, w322, g2);
and (w324, w323, w313);
or (w325, w324, w285);
and (w326, w325, g6);
or (w327, w326, w226);
or (w328, w327, w145);
or (w329, w328, w70);
or (w330, w329, w131);
and (w331, w131, w47);
and (w332, g7, g3);
and (w333, w332, w103);
or (w334, g7, g3);
or (w335, w334, w301);
and (w336, w335, w51);
or (w337, w336, w333);
or (w338, g9, g8);
and (w339, w338, w66);
or (w340, w339, w3);
and (w341, g7, g3);
and (w342, w341, w103);
or (w343, g7, g3);
or (w344, w343, w301);
and (w345, w344, w51);
or (w346, w345, w342);
and (w347, w346, w337);
and (w348, w347, w340);
or (w349, w348, w331);
and (w350, w333, g7);
and (w351, w350, g3);
and (w352, w351, w103);
and (w353, w352, w340);
or (w354, w353, w331);
or (w355, w340, w331);
or (w356, g7, g3);
and (w357, w355, w356);
or (w358, w357, w301);
and (w359, w358, w51);
or (w360, w359, w354);
and (w361, w360, w349);
and (w362, w361, w340);
or (w363, w362, w331);
and (w364, w363, w330);
or (w365, w131, w340);
and (w366, w365, g7);
and (w367, w366, g3);
and (w368, w367, w103);
or (w369, w51, w368);
and (w370, w369, w356);
or (w371, w370, w301);
and (w372, w371, w51);
or (w373, w372, w368);
or (w374, w131, w340);
and (w375, w374, w373);
and (w376, w375, w131);
or (w377, w376, w340);
and (w378, w377, w373);
and (w379, w364, w378);
and (w380, w3, w379);
and (w381, w340, w379);
or (w382, w131, w381);
and (w383, w379, w382);
and (w384, w379, w382);
and (w385, w384, w383);
or (w386, g1, g5);
or (w387, w381, g1);
or (w388, w387, g1);
or (w389, w388, g5);
and (w390, w389, w386);
or (w391, w381, g1);
or (w392, w391, g1);
or (w393, w392, g5);
or (w394, w381, g9);
or (w395, w394, g8);
and (w396, w395, g9);
and (w397, w396, g8);
or (w398, w397, w380);
and (w399, w382, w379);
or (w400, w390, w381);
or (w401, w400, w398);
or (w402, w401, w398);
or (w403, w402, w381);
or (w404, w403, g2);
or (w405, w404, g2);
or (w406, w390, w381);
or (w407, w406, w398);
or (w408, w407, w398);
or (w409, w408, w381);
or (w410, w409, g2);
or (w411, w410, g2);
and (w412, w411, w405);
or (w413, w412, w381);
or (w414, w398, w381);
or (w415, w414, g1);
or (w416, w415, g1);
and (w417, w416, w393);
or (w418, w417, w413);
and (w419, w418, w382);
and (w420, w419, w379);
and (w421, w420, w364);
and (w422, w421, w378);
or (w423, w422, g6);
or (w424, w423, g6);
and (w425, w424, w385);
and (w426, w382, w379);
and (w427, w426, w364);
and (w428, w427, w378);
and (w429, w428, w390);
or (w430, w429, w381);
and (w431, w430, w379);
or (w432, w431, w381);
and (w433, w432, w382);
or (w434, w433, w398);
or (w435, w434, w398);
or (w436, w435, w381);
or (w437, w436, g2);
or (w438, w437, g2);
or (w439, w438, g6);
or (w440, w439, g6);
and (w441, w440, w425);
or (w442, w398, w381);
or (w443, w442, g1);
or (w444, w443, g1);
or (w445, w444, g5);
or (w446, w445, g5);
or (w447, w381, w398);
or (w448, w447, g1);
or (w449, w448, g1);
or (w450, w449, g5);
or (w451, w450, g5);
and (w452, w451, w446);
and (w453, w452, w382);
and (w454, w453, w379);
and (w455, w454, w364);
and (w456, w455, w378);
and (w457, w456, w379);
or (w458, w457, w381);
and (w459, w458, w382);
or (w460, w459, w398);
or (w461, w460, w398);
or (w462, w461, w381);
or (w463, w462, g2);
or (w464, w463, g2);
and (w465, w464, w441);
or (w466, w465, g6);
or (w467, w466, g6);
and (w468, w467, w425);
or (w469, w37, w398);
or (w470, w469, w19);
or (w471, w470, w16);
or (w472, w471, w381);
or (w473, w472, w398);
or (w474, w473, w398);
or (w475, w474, w381);
or (w476, w475, g2);
or (w477, w476, g2);
or (w478, w37, w398);
or (w479, w478, w19);
or (w480, w479, w16);
or (w481, w480, w381);
or (w482, w481, w398);
or (w483, w482, w398);
or (w484, w483, w381);
or (w485, w484, g2);
or (w486, w485, g2);
and (w487, w486, w477);
or (w488, w487, w468);
or (w489, w488, g6);
or (w490, w489, g6);
and (w491, w490, w425);
or (w492, w491, w398);
or (w493, w492, w381);
or (w494, w493, w54);
or (w495, w494, g3);
or (w496, w495, g3);
or (w497, w37, w398);
or (w498, w497, w19);
or (w499, w498, w16);
or (w500, w499, w381);
or (w501, w500, w398);
or (w502, w501, w398);
or (w503, w502, w381);
or (w504, w503, g2);
or (w505, w504, g2);
and (w506, w505, w477);
or (w507, w506, g6);
or (w508, w507, g6);
or (w509, w508, w468);
and (w510, w509, w425);
or (w511, w510, w398);
or (w512, w511, w398);
or (w513, w512, w381);
or (w514, w513, w381);
or (w515, w514, g3);
or (w516, w515, g3);
and (w517, w516, w496);
and (w518, w517, w399);
or (w519, w518, g7);
or (w520, w519, g7);
and (w521, g7, w520);
and (w522, g7, w520);
and (w523, w379, w382);
and (w524, w523, w364);
and (w525, w524, w378);
and (w526, w525, w390);
and (w527, w526, w379);
and (w528, w527, w382);
and (w529, w528, w379);
and (w530, w529, w382);
or (w531, w530, w398);
or (w532, w531, w398);
or (w533, w532, w398);
or (w534, w533, w381);
or (w535, w534, w381);
and (w536, w535, w520);
and (w537, w536, w520);
and (w538, w537, w520);
or (w539, w538, w522);
or (w540, w539, w381);
and (w541, w540, w103);
or (w542, w541, w521);
and (w543, w542, g3);
or (w544, w543, w301);
and (w545, w468, w382);
or (w546, w545, w398);
or (w547, w546, w398);
and (w548, w547, w520);
or (w549, w548, w522);
or (w550, w549, w381);
and (w551, w550, w379);
or (w552, w551, w381);
or (w553, w552, g3);
and (w554, w553, w520);
or (w555, w554, w521);
and (w556, w555, g3);
and (w557, w556, w520);
or (w558, w557, w521);
and (w559, w558, w356);
or (w560, w381, w544);
or (w561, w560, g6);
and (w562, w561, g6);
or (w563, w562, w398);
or (w564, w563, w381);
or (w565, w564, w559);
or (w566, w381, w398);
or (w567, w566, g1);
or (w568, w567, g1);
or (w569, w568, g5);
or (w570, w569, g5);
and (w571, w570, w446);
and (w572, w571, w382);
and (w573, w572, w379);
and (w574, w573, w364);
and (w575, w574, w378);
and (w576, w575, w379);
or (w577, w576, w381);
and (w578, w577, w382);
or (w579, w578, w398);
or (w580, w579, g6);
and (w581, w580, g6);
or (w582, w581, w565);
or (w583, w582, w398);
or (w584, w583, w381);
or (w585, w584, g2);
or (w586, w585, g2);
and (w587, w586, w379);
and (w588, w587, w382);
or (w589, w588, w398);
or (w590, w589, w398);
or (w591, w590, w381);
and (w592, w591, w520);
and (w593, w592, w520);
and (w594, w593, w520);
or (w595, w594, w522);
or (w596, w595, w381);
and (w597, w596, w103);
or (w598, w597, w521);
and (w599, w598, g3);
or (w600, w599, w301);
or (w601, w600, w559);
or (w602, w381, w398);
or (w603, w602, g1);
or (w604, w603, g1);
or (w605, w604, g5);
or (w606, w605, g5);
and (w607, w606, w446);
and (w608, w607, w382);
and (w609, w608, w379);
and (w610, w609, w364);
and (w611, w610, w378);
and (w612, w611, w379);
or (w613, w612, w381);
and (w614, w613, w382);
or (w615, w614, w398);
or (w616, w615, g6);
and (w617, w616, g6);
or (w618, w617, w398);
or (w619, w618, w381);
or (w620, w619, g2);
or (w621, w620, g2);
and (w622, w621, w601);
and (w623, w622, w379);
and (w624, w623, w382);
or (w625, w624, w398);
or (w626, w625, w398);
or (w627, w626, w381);
and (w628, w627, w520);
and (w629, w628, w520);
and (w630, w629, w520);
or (w631, w630, w522);
or (w632, w631, w381);
and (w633, w632, w103);
or (w634, w633, w521);
and (w635, w634, g3);
or (w636, w635, w301);
or (w637, w636, w559);
or (w638, w381, w398);
or (w639, w638, g1);
or (w640, w639, g1);
or (w641, w640, g5);
or (w642, w641, g5);
and (w643, w642, w446);
and (w644, w643, w382);
and (w645, w644, w379);
and (w646, w645, w364);
and (w647, w646, w378);
and (w648, w647, w379);
or (w649, w648, w381);
and (w650, w649, w382);
or (w651, w650, w398);
or (w652, w651, g6);
and (w653, w652, g6);
or (w654, w653, w637);
or (w655, w654, w398);
or (w656, w655, w381);
or (w657, w656, g2);
or (w658, w657, g2);
and (w659, w658, w601);
and (w660, w659, w379);
and (w661, w660, w382);
or (w662, w661, w398);
or (w663, w662, w398);
or (w664, w663, w381);
and (w665, w664, w520);
and (w666, w665, w520);
and (w667, w666, w520);
or (w668, w667, w522);
or (w669, w668, w381);
and (w670, w669, w103);
or (w671, w670, w521);
and (w672, w671, g3);
or (w673, w672, w301);
or (w674, w673, w559);
or (w675, w674, w398);
or (w676, w675, w381);
or (w677, w676, g1);
or (w678, w677, g1);
and (w679, g1, w678);
and (w680, g1, w678);
or (w681, w679, w381);
or (w682, w680, w398);
or (w683, w681, w674);
or (w684, w682, w683);
endmodule