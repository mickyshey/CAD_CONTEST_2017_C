module patch (w43, a, b, c, g1);
input a, b, c, g1;
output w43;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43;
not(w0, g1);
or (w1, w0, a);
not(w2, g1);
or (w3, w2, b);
not(w4, a);
or (w5, g1, w4);
not(w6, b);
or (w7, w5, w6);
not(w8, b);
not(w9, c);
not(w10, c);
not(w11, a);
or (w12, w11, c);
not(w13, a);
not(w14, b);
not(w15, c);
not(w16, b);
or (w17, w15, w16);
or (w18, g1, b);
and (w19, w18, w3);
and (w20, g1, w1);
and (w21, w20, w12);
and (w22, w21, w17);
or (w23, w22, w8);
and (w24, w23, w19);
or (w25, w24, w10);
or (w26, w25, w9);
or (w27, w26, w13);
or (w28, w27, b);
or (w29, c, w24);
or (w30, w29, a);
and (w31, w30, w7);
or (w32, w31, w14);
or (w33, w32, w8);
and (w34, w33, w28);
and (w35, w1, w34);
and (w36, w3, w34);
and (w37, w35, w36);
and (w38, w37, w35);
and (w39, w37, w35);
and (w40, w38, w36);
and (w41, w39, w34);
and (w42, w41, w40);
and (w43, w42, w38);
endmodule