module patch (1'b0, 
input 
output 1'b0;
wire 
endmodule
