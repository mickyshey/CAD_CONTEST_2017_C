module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 ;
output g11 , g12 , g13 , g14 , g15 , g16 ;
wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 ;
wire t_0 , w5 , w6 , w7 , w63 , w64 , w360 , w18 , w19 , w46 , w47 , w332 , w48 , w49 , w21 , w22 , w146 , w333 , w74 , w75 , w76 , w334 , w60 , w335 , w28 , w29 , w99 , w69 , w26 , w27 , w98 , w100 , w77 , w78 , w79 , w101 , w102 , w103 , w14 , w15 , w16 , w95 , w96 , w30 , w31 , w32 , w72 , w73 , w93 , w25 , w70 , w71 , w92 , w94 , w97 , w104 , w336 , w259 , w260 , w59 , w261 , w262 , w50 , w51 , w52 , w61 , w250 , w13 , w251 , w39 , w40 , w41 , w53 , w54 , w55 , w179 , w180 , w181 , w35 , w36 , w111 , w44 , w112 , w87 , w113 , w83 , w114 , w115 , w82 , w37 , w38 , w106 , w34 , w84 , w105 , w107 , w108 , w109 , w110 , w116 , w174 , w175 , w176 , w85 , w42 , w119 , w120 , w177 , w43 , w86 , w117 , w118 , w178 , w182 , w183 , w184 , w185 , w186 , w187 , w252 , w253 , w233 , w234 , w224 , w225 , w226 , w227 , w207 , w208 , w209 , w210 , w45 , w88 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w159 , w160 , w161 , w162 , w163 , w164 , w147 , w148 , w149 , w56 , w57 , w58 , w150 , w151 , w152 , w153 , w133 , w134 , w135 , w136 , w121 , w122 , w123 , w124 , w125 , w126 , w127 , w128 , w129 , w130 , w131 , w65 , w62 , w90 , w89 , w91 , w132 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w154 , w155 , w156 , w157 , w158 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w203 , w204 , w205 , w206 , w211 , w212 , w213 , w214 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w228 , w229 , w230 , w231 , w232 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w254 , w255 , w256 , w257 , w258 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w337 , w338 , w339 , w340 , w341 , w342 , w302 , w303 , w304 , w305 , w306 , w284 , w285 , w286 , w287 , w288 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w307 , w308 , w309 , w310 , w311 , w343 , w344 , w345 , w346 , w347 , w3 , w4 , w348 , w349 , w350 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w1 , w2 , w328 , w329 , w330 , w331 , w351 , w352 , w361 , w0 , w66 , w67 , w358 , w359 , w362 , w963 , w964 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w81 , w737 , w738 , w33 , w739 , w740 , w432 , w431 , w433 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w80 , w717 , w718 , w719 , w24 , w720 , w721 , w722 , w434 , w435 , w436 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w700 , w701 , w702 , w723 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w654 , w675 , w676 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w451 , w452 , w453 , w454 , w455 , w456 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w650 , w651 , w652 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w12 , w624 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w8 , w9 , w10 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w353 , w354 , w355 , w356 , w357 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w481 , w482 , w483 , w484 , w485 , w526 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w11 , w569 , w570 , w582 , w583 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w511 , w512 , w513 , w514 , w515 , w516 , w545 , w546 , w547 , w548 , w549 , w550 , w584 , w585 , w586 , w587 , w588 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w653 , w677 , w678 , w679 , w680 , w681 , w682 , w724 , w725 , w726 , w727 , w728 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w68 , w760 , w23 , w761 , w762 , w757 , w758 , w759 , w763 , w764 , w965 , w966 , w967 , w20 , w765 , w792 , w793 , w17 , w794 , w795 , w796 , w968 , w902 , w903 , w904 , w905 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w843 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w842 , w862 , w863 , w864 , w865 , w866 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w867 , w898 , w899 , w900 , w901 , w921 , w922 , w923 , w924 , w925 , w926 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1013 , w1014 , w1015 , w1016 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w927 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w928 , w929 , w930 , w931 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w996 , w997 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1062 , w1063 , w1067 , w1073 , w1065 , w1072 , w1076 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1068 , w1069 , w1097 , w1098 , w1071 , w1099 , w1100 , w1070 , w1101 , w1075 , w1074 , w1077 , w1102 , w1064 , w1103 , w1066 , w1104 , w1107 , w1108 , w1061 , w1110 , w1112 , w1113 , w1105 , w1106 , w1060 , w1109 , w1114 , w1111 , w1115;
buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( g11 , n12  );
buf ( g12 , n13  );
buf ( g13 , n14  );
buf ( g14 , n15  );
buf ( g15 , n16  );
buf ( g16 , n17  );
buf ( n12 , n40 );
buf ( n13 , n65 );
buf ( n14 , n70 );
buf ( n15 , n44 );
buf ( n16 , n54 );
buf ( n17 , n60 );
xnor ( n20 , n9 , n10 );
not ( n21 , n3 );
not ( n22 , n7 );
or ( n23 , n21 , n22 );
nor ( n24 , n3 , n7 );
not ( n25 , n24 );
nand ( n26 , n4 , n8 );
not ( n27 , n26 );
nand ( n28 , n25 , n27 );
nand ( n29 , n23 , n28 );
not ( n30 , n2 );
and ( n31 , n6 , n30 );
not ( n32 , n6 );
and ( n33 , n32 , n2 );
nor ( n34 , n31 , n33 );
and ( n35 , n29 , n34 );
nor ( n36 , n35 , t_0 );
or ( n37 , n20 , n36 );
not ( n38 , n20 );
or ( n39 , n30 , n38 );
nand ( n40 , n37 , n39 );
or ( n41 , n38 , n36 );
not ( n42 , n6 );
or ( n43 , n42 , n20 );
nand ( n44 , n41 , n43 );
not ( n45 , n7 );
not ( n46 , n38 );
or ( n47 , n45 , n46 );
xor ( n48 , n3 , n7 );
and ( n49 , n48 , n26 );
not ( n50 , n48 );
and ( n51 , n50 , n27 );
nor ( n52 , n49 , n51 );
or ( n53 , n52 , n38 );
nand ( n54 , n47 , n53 );
not ( n55 , n8 );
not ( n56 , n38 );
or ( n57 , n55 , n56 );
xnor ( n58 , n4 , n8 );
or ( n59 , n58 , n38 );
nand ( n60 , n57 , n59 );
not ( n61 , n3 );
not ( n62 , n20 );
or ( n63 , n61 , n62 );
or ( n64 , n20 , n52 );
nand ( n65 , n63 , n64 );
not ( n66 , n4 );
not ( n67 , n20 );
or ( n68 , n66 , n67 );
or ( n69 , n58 , n20 );
nand ( n70 , n68 , n69 );
buf ( t_0, w1115 );
not(w5, g9);
not(w6, g8);
or (w7, w5, w6);
not(w63, g9);
or (w64, w63, g8);
and (w360, w7, w64);
not(w18, g5);
or (w19, g1, w18);
not(w46, g5);
or (w47, g1, w46);
or (w332, w19, w47);
not(w48, g1);
or (w49, w48, g5);
not(w21, g1);
or (w22, w21, g5);
or (w146, w49, w22);
and (w333, w332, w146);
not(w74, g2);
not(w75, g6);
or (w76, w74, w75);
and (w334, w333, w76);
not(w60, g6);
or (w335, w334, w60);
not(w28, g2);
or (w29, w28, g6);
and (w99, w76, w29);
or (w69, g2, g6);
not(w26, g6);
or (w27, g2, w26);
and (w98, w69, w27);
and (w100, w99, w98);
not(w77, g3);
not(w78, g7);
or (w79, w77, w78);
or (w101, w100, w79);
and (w102, w101, g7);
and (w103, w102, g3);
not(w14, g3);
not(w15, g7);
or (w16, w14, w15);
and (w95, w16, g7);
and (w96, w95, g3);
not(w30, g2);
not(w31, g6);
or (w32, w30, w31);
not(w72, g2);
or (w73, w72, g6);
and (w93, w32, w73);
or (w25, g2, g6);
not(w70, g6);
or (w71, g2, w70);
and (w92, w25, w71);
and (w94, w93, w92);
or (w97, w96, w94);
or (w104, w103, w97);
or (w336, w335, w104);
or (w259, w19, w47);
or (w260, w259, w104);
not(w59, g2);
or (w261, w260, w59);
and (w262, w261, w69);
not(w50, g1);
not(w51, g5);
or (w52, w50, w51);
or (w61, g2, g6);
or (w250, w52, w61);
or (w13, g2, g6);
or (w251, w250, w13);
not(w39, g3);
not(w40, g7);
or (w41, w39, w40);
not(w53, g3);
not(w54, g7);
or (w55, w53, w54);
or (w179, w41, w55);
or (w180, w179, w16);
or (w181, w180, w79);
not(w35, g7);
or (w36, g3, w35);
or (w111, w36, g3);
not(w44, g7);
or (w112, w111, w44);
not(w87, g7);
or (w113, w112, w87);
not(w83, g7);
or (w114, w113, w83);
and (w115, w114, w16);
not(w82, g3);
not(w37, g3);
or (w38, w37, g7);
or (w106, w82, w38);
or (w34, g3, g7);
or (w84, g3, g7);
or (w105, w34, w84);
and (w107, w106, w105);
or (w108, w107, g7);
or (w109, w108, g7);
or (w110, w109, g7);
and (w116, w115, w110);
or (w174, w116, g3);
or (w175, w174, g3);
or (w176, w175, w94);
not(w85, g5);
not(w42, g5);
or (w119, w85, w42);
and (w120, w119, g5);
or (w177, w176, w120);
not(w43, g6);
not(w86, g6);
or (w117, w43, w86);
and (w118, w117, g6);
or (w178, w177, w118);
and (w182, w181, w178);
or (w183, w182, w94);
or (w184, w183, w44);
or (w185, w184, w87);
or (w186, w185, w120);
or (w187, w186, w118);
or (w252, w251, w187);
and (w253, w252, w73);
or (w233, w52, w29);
and (w234, w233, w69);
or (w224, w52, w187);
and (w225, w224, w73);
or (w226, w225, g3);
or (w227, w226, g3);
or (w207, w146, w104);
or (w208, w207, w41);
or (w209, w208, w55);
or (w210, w209, w79);
or (w45, g1, g5);
and (w88, w49, g1);
or (w195, w45, w88);
or (w196, w195, w36);
or (w197, w196, g3);
or (w198, w197, g3);
or (w199, w198, g3);
or (w200, w199, w44);
or (w201, w200, w87);
or (w202, w201, w83);
and (w159, w52, w45);
or (w160, w159, w110);
or (w161, w160, w27);
or (w162, w161, g2);
or (w163, w162, g2);
and (w164, w163, w76);
or (w147, w19, w47);
and (w148, w147, w146);
or (w149, w148, w110);
not(w56, g2);
not(w57, g6);
or (w58, w56, w57);
or (w150, w149, w58);
or (w151, w150, w104);
and (w152, w151, w71);
or (w153, w152, w60);
and (w133, w52, w45);
or (w134, w133, w110);
or (w135, w134, w29);
and (w136, w135, w69);
and (w121, w52, w45);
or (w122, w121, w110);
or (w123, w122, w104);
and (w124, w123, w73);
or (w125, w124, g6);
or (w126, w125, g6);
or (w127, w126, g7);
or (w128, w127, g7);
or (w129, w128, g7);
or (w130, w129, w120);
or (w131, w130, w118);
not(w65, g9);
not(w62, g8);
or (w90, w65, w62);
or (w89, g9, g8);
and (w91, w90, w89);
and (w132, w131, w91);
or (w137, w136, w132);
or (w138, w137, g6);
or (w139, w138, g6);
or (w140, w139, g7);
or (w141, w140, g7);
or (w142, w141, g7);
or (w143, w142, w120);
or (w144, w143, w118);
and (w145, w144, w91);
and (w154, w153, w145);
or (w155, w154, g7);
or (w156, w155, w120);
or (w157, w156, w118);
and (w158, w157, w91);
or (w165, w164, w158);
and (w166, w165, w145);
or (w167, w166, g7);
or (w168, w167, g7);
or (w169, w168, g7);
or (w170, w169, w120);
or (w171, w170, w118);
and (w172, w171, w91);
and (w173, w172, w91);
and (w203, w202, w173);
or (w204, w203, w120);
or (w205, w204, w118);
and (w206, w205, w91);
and (w211, w210, w206);
or (w212, w211, w59);
or (w213, w212, w29);
and (w214, w213, w69);
or (w188, w45, w187);
or (w189, w188, w61);
or (w190, w189, w13);
and (w191, w190, w73);
or (w192, w191, g6);
and (w193, w192, w173);
and (w194, w193, w91);
or (w215, w214, w194);
or (w216, w215, g6);
or (w217, w216, g6);
or (w218, w217, w44);
or (w219, w218, w87);
and (w220, w219, w173);
or (w221, w220, w120);
or (w222, w221, w118);
and (w223, w222, w91);
and (w228, w227, w223);
or (w229, w228, g6);
or (w230, w229, g6);
and (w231, w230, w173);
and (w232, w231, w91);
or (w235, w234, w232);
or (w236, w235, w36);
or (w237, w236, g3);
or (w238, w237, g3);
or (w239, w238, g3);
and (w240, w239, w223);
or (w241, w240, g6);
or (w242, w241, g6);
or (w243, w242, w44);
or (w244, w243, w87);
or (w245, w244, w83);
and (w246, w245, w173);
or (w247, w246, w120);
or (w248, w247, w118);
and (w249, w248, w91);
and (w254, w253, w249);
and (w255, w254, w223);
or (w256, w255, g6);
and (w257, w256, w173);
and (w258, w257, w91);
or (w263, w262, w258);
or (w264, w263, w41);
or (w265, w264, w55);
or (w266, w265, w79);
and (w267, w266, w249);
and (w268, w267, w223);
or (w269, w268, w44);
or (w270, w269, w87);
and (w271, w270, w173);
or (w272, w271, w120);
or (w273, w272, w118);
and (w274, w273, w91);
and (w337, w336, w274);
or (w338, w337, w41);
or (w339, w338, w55);
or (w340, w339, w79);
or (w341, w340, w44);
or (w342, w341, w87);
or (w302, w19, w47);
and (w303, w302, w146);
and (w304, w303, w71);
or (w305, w304, w187);
or (w306, w305, w55);
and (w284, w52, w206);
or (w285, w284, w27);
or (w286, w285, g2);
or (w287, w286, g2);
and (w288, w287, w76);
or (w275, w19, w47);
and (w276, w275, w146);
or (w277, w276, w58);
and (w278, w277, w71);
or (w279, w278, w187);
or (w280, w279, w60);
and (w281, w280, w274);
and (w282, w281, w173);
and (w283, w282, w91);
or (w289, w288, w283);
or (w290, w289, w36);
or (w291, w290, g3);
or (w292, w291, g3);
or (w293, w292, g3);
and (w294, w293, w274);
or (w295, w294, w44);
or (w296, w295, w87);
or (w297, w296, w83);
and (w298, w297, w173);
or (w299, w298, w120);
or (w300, w299, w118);
and (w301, w300, w91);
and (w307, w306, w301);
or (w308, w307, w60);
and (w309, w308, w274);
and (w310, w309, w173);
and (w311, w310, w91);
or (w343, w342, w311);
and (w344, w343, w301);
and (w345, w344, w173);
or (w346, w345, w120);
or (w347, w346, w118);
not(w3, g8);
or (w4, g9, w3);
or (w348, w347, w4);
and (w349, w348, g8);
and (w350, w349, w65);
or (w312, w19, w47);
and (w313, w312, w146);
or (w314, w313, w104);
and (w315, w314, w76);
or (w316, w315, w311);
or (w317, w316, w41);
or (w318, w317, w55);
or (w319, w318, w79);
and (w320, w319, w301);
or (w321, w320, w60);
and (w322, w321, w274);
or (w323, w322, w44);
or (w324, w323, w87);
and (w325, w324, w173);
or (w326, w325, w120);
or (w327, w326, w118);
not(w1, g9);
or (w2, w1, g8);
or (w328, w327, w2);
and (w329, w328, w62);
and (w330, w329, g9);
and (w331, w330, w91);
or (w351, w350, w331);
and (w352, w351, w91);
or (w361, w360, w352);
or (w0, g9, g8);
not(w66, g8);
or (w67, g9, w66);
and (w358, w0, w67);
or (w359, w358, w352);
and (w362, w361, w359);
or (w963, w362, w352);
or (w964, w963, w19);
or (w729, g5, w362);
or (w730, w729, w352);
or (w731, w730, w352);
or (w732, w731, w362);
or (w733, w732, w104);
or (w734, w733, w41);
or (w735, w734, w55);
or (w736, w735, w79);
not(w81, g3);
or (w737, w736, w81);
or (w738, w737, w352);
not(w33, g3);
or (w739, w738, w33);
or (w740, w739, w362);
or (w432, w64, w352);
or (w431, w67, w352);
and (w433, w432, w431);
and (w741, w740, w433);
and (w742, w741, w433);
and (w743, w742, w433);
or (w744, w743, w352);
or (w745, w744, w362);
or (w746, w745, g2);
or (w747, w746, g2);
and (w748, w747, w76);
or (w749, w748, w60);
or (w703, g5, g6);
or (w704, w703, w352);
or (w705, w704, w362);
or (w706, w705, w104);
or (w707, w706, w41);
or (w708, w707, w55);
or (w709, w708, w79);
or (w710, w709, w81);
or (w711, w710, w352);
or (w712, w711, w33);
or (w713, w712, w362);
and (w714, w713, w433);
and (w715, w714, w433);
and (w716, w715, w433);
not(w80, g2);
or (w717, w716, w80);
or (w718, w717, w352);
or (w719, w718, w59);
not(w24, g2);
or (w720, w719, w24);
or (w721, w720, w362);
and (w722, w721, w69);
and (w434, w433, w45);
and (w435, w434, w433);
and (w436, w435, w45);
and (w693, w433, w436);
and (w694, w693, w433);
and (w695, w694, w433);
and (w696, w695, w433);
and (w697, w696, w433);
and (w698, w697, w433);
and (w699, w698, w76);
and (w683, w433, w436);
and (w684, w683, w433);
and (w685, w684, w433);
and (w686, w685, w433);
and (w687, w686, w433);
and (w688, w687, w433);
and (w689, w688, w433);
and (w690, w689, w69);
and (w691, w690, w433);
and (w692, w691, w45);
and (w700, w699, w692);
and (w701, w700, w433);
and (w702, w701, w45);
and (w723, w722, w702);
or (w655, w362, w352);
or (w656, w655, w362);
or (w657, w656, w352);
or (w658, w657, w362);
or (w659, w658, w352);
or (w660, w659, w36);
or (w661, w660, g3);
or (w662, w661, g3);
or (w663, w662, g3);
or (w664, w663, g3);
and (w665, w664, w55);
or (w397, w362, w352);
or (w398, w397, w352);
or (w399, w398, w41);
or (w400, w399, w16);
or (w401, w400, w79);
or (w402, w401, w81);
or (w403, w402, w352);
or (w404, w403, w33);
or (w405, w404, w362);
and (w406, w405, g3);
or (w407, w406, w94);
or (w666, w665, w407);
or (w667, w666, g5);
or (w668, w667, w58);
or (w669, w668, w80);
or (w670, w669, w352);
or (w671, w670, w24);
or (w672, w671, w362);
and (w673, w672, w71);
or (w674, w673, w60);
and (w654, w433, w73);
and (w675, w674, w654);
or (w676, w675, w83);
or (w444, w362, w38);
or (w445, w444, w81);
or (w446, w445, w352);
or (w447, w446, w33);
or (w448, w447, w362);
and (w449, w448, w84);
or (w450, w449, w352);
or (w437, w362, w105);
or (w438, w437, w34);
or (w439, w438, g3);
or (w440, w439, g3);
and (w441, w440, w82);
or (w442, w441, w352);
or (w443, w442, g7);
or (w451, w450, w443);
or (w452, w451, w362);
or (w453, w452, w352);
or (w454, w453, g7);
or (w455, w454, g7);
or (w456, w455, w94);
or (w642, g5, w456);
or (w643, w642, w58);
or (w644, w643, w80);
or (w645, w644, w352);
or (w646, w645, w24);
or (w647, w646, w362);
and (w648, w647, w71);
or (w649, w648, w60);
and (w632, w433, w436);
and (w633, w632, w433);
and (w634, w633, w433);
and (w635, w634, w433);
and (w636, w635, w433);
and (w637, w636, w433);
and (w638, w637, w433);
and (w639, w638, w73);
and (w640, w639, w433);
and (w641, w640, w45);
and (w650, w649, w641);
or (w651, w650, w22);
and (w652, w651, w45);
or (w602, g5, w362);
or (w603, w602, w352);
or (w604, w603, w362);
or (w605, w604, w352);
or (w606, w605, w362);
or (w607, w606, w352);
or (w608, w607, w36);
or (w609, w608, g3);
or (w610, w609, g3);
or (w611, w610, g3);
or (w612, w611, g3);
and (w613, w612, w55);
or (w589, w362, w352);
or (w590, w589, w352);
or (w591, w590, w362);
or (w592, w591, w104);
or (w593, w592, w352);
or (w594, w593, w41);
or (w595, w594, w16);
or (w596, w595, w79);
or (w597, w596, w81);
or (w598, w597, w352);
or (w599, w598, w33);
or (w600, w599, w362);
and (w601, w600, g3);
or (w614, w613, w601);
or (w615, w614, w352);
or (w616, w615, w362);
or (w617, w616, w27);
or (w618, w617, g2);
or (w619, w618, g2);
or (w620, w619, g2);
or (w621, w620, g2);
and (w622, w621, w76);
or (w623, w622, w60);
not(w12, g6);
or (w624, w623, w12);
or (w517, g5, w362);
or (w518, w517, w80);
or (w519, w518, w352);
or (w520, w519, w29);
or (w521, w520, w24);
or (w522, w521, w362);
and (w523, w522, w69);
or (w524, w523, g6);
or (w525, w524, g6);
or (w457, w362, w352);
or (w458, w457, w362);
or (w459, w458, w352);
or (w460, w459, w362);
or (w461, w460, w36);
or (w462, w461, g3);
or (w463, w462, g3);
or (w464, w463, g3);
or (w465, w464, g3);
or (w466, w465, w352);
and (w467, w466, w55);
or (w468, w467, w407);
or (w469, w468, w83);
and (w470, w469, w456);
or (w471, w470, w352);
or (w472, w471, w362);
or (w473, w472, w58);
not(w8, g2);
not(w9, g6);
or (w10, w8, w9);
or (w474, w473, w10);
or (w475, w474, w80);
or (w476, w475, w352);
or (w477, w476, w24);
or (w478, w477, w362);
and (w479, w478, w71);
or (w480, w479, w60);
or (w408, g6, w362);
or (w409, w408, w352);
or (w410, w409, w362);
or (w411, w410, w352);
or (w412, w411, w36);
or (w413, w412, g3);
or (w414, w413, g3);
or (w415, w414, g3);
or (w416, w415, g3);
and (w417, w416, w55);
or (w418, w417, w407);
or (w419, w418, w83);
or (w353, g5, w352);
or (w354, w353, g2);
and (w355, w354, w73);
or (w356, w355, g6);
or (w357, w356, g6);
or (w379, w357, w352);
or (w380, w379, w362);
or (w381, w380, w38);
or (w382, w381, w82);
or (w383, w382, w81);
or (w384, w383, w352);
or (w385, w384, w33);
or (w386, w385, w362);
or (w363, w352, w362);
or (w364, w363, w357);
or (w365, w364, w105);
or (w366, w365, w34);
or (w367, w366, w84);
or (w368, w367, g3);
or (w369, w368, g3);
or (w370, w369, g7);
or (w371, w370, g7);
or (w372, w371, g7);
or (w373, w372, w362);
or (w374, w373, w13);
or (w375, w374, g2);
and (w376, w375, w73);
or (w377, w376, w94);
or (w378, w377, g6);
and (w387, w386, w378);
or (w388, w387, g7);
or (w389, w388, g7);
or (w390, w389, g7);
or (w391, w390, w362);
or (w392, w391, w13);
or (w393, w392, g2);
and (w394, w393, w73);
or (w395, w394, w94);
or (w396, w395, g6);
and (w420, w419, w396);
or (w421, w420, g5);
or (w422, w421, w352);
or (w423, w422, w362);
or (w424, w423, w61);
or (w425, w424, w13);
or (w426, w425, g2);
or (w427, w426, g2);
and (w428, w427, w73);
or (w429, w428, w94);
or (w430, w429, g6);
and (w481, w480, w430);
or (w482, w481, w94);
or (w483, w482, g1);
and (w484, w483, w49);
or (w485, w484, g5);
or (w526, w525, w485);
or (w571, w526, w352);
or (w572, w571, w362);
or (w573, w572, w352);
or (w574, w573, w362);
or (w575, w574, w352);
or (w576, w575, w36);
or (w577, w576, g3);
or (w578, w577, g3);
or (w579, w578, g3);
or (w580, w579, g3);
and (w581, w580, w55);
or (w551, w362, g6);
or (w552, w551, w352);
or (w553, w552, w362);
or (w554, w553, w104);
or (w555, w554, w352);
or (w556, w555, w41);
or (w557, w556, w16);
or (w558, w557, w79);
or (w559, w558, w81);
or (w560, w559, w352);
or (w561, w560, w33);
or (w562, w561, w362);
and (w563, w562, g3);
or (w564, w563, w80);
or (w565, w564, w352);
or (w566, w565, w59);
or (w567, w566, w24);
or (w568, w567, w362);
not(w11, g2);
or (w569, w568, w11);
and (w570, w569, w69);
or (w582, w581, w570);
or (w583, w582, w83);
or (w527, g5, w362);
or (w528, w527, w352);
or (w529, w528, w362);
or (w530, w529, w27);
or (w531, w530, g2);
or (w532, w531, g2);
or (w533, w532, g2);
or (w534, w533, g2);
and (w535, w534, w76);
and (w536, w535, w526);
or (w537, w536, w362);
or (w538, w537, w38);
or (w539, w538, w81);
or (w540, w539, w352);
or (w541, w540, w33);
or (w542, w541, w362);
and (w543, w542, w84);
or (w544, w543, w352);
or (w501, w443, g5);
or (w502, w501, w362);
or (w503, w502, w352);
or (w504, w503, w362);
or (w505, w504, w27);
or (w506, w505, g2);
or (w507, w506, g2);
or (w508, w507, g2);
or (w509, w508, g2);
and (w510, w509, w76);
or (w486, w443, g5);
or (w487, w486, w362);
or (w488, w487, w80);
or (w489, w488, w352);
or (w490, w489, w29);
or (w491, w490, w24);
or (w492, w491, w362);
and (w493, w492, w69);
or (w494, w493, g6);
or (w495, w494, g6);
or (w496, w495, w352);
or (w497, w496, g7);
or (w498, w497, g7);
or (w499, w498, g7);
or (w500, w499, w485);
and (w511, w510, w500);
or (w512, w511, w352);
or (w513, w512, g7);
or (w514, w513, g7);
or (w515, w514, g7);
or (w516, w515, w485);
or (w545, w544, w516);
or (w546, w545, w352);
or (w547, w546, g7);
or (w548, w547, g7);
or (w549, w548, g7);
or (w550, w549, w485);
and (w584, w583, w550);
or (w585, w584, w485);
or (w586, w585, g1);
and (w587, w586, w49);
or (w588, w587, g5);
and (w625, w624, w588);
or (w626, w625, w83);
and (w627, w626, w550);
or (w628, w627, w485);
or (w629, w628, g1);
and (w630, w629, w49);
or (w631, w630, g5);
or (w653, w652, w631);
and (w677, w676, w653);
or (w678, w677, w94);
and (w679, w678, w433);
or (w680, w679, w22);
and (w681, w680, w45);
or (w682, w681, w631);
or (w724, w723, w682);
and (w725, w724, w433);
or (w726, w725, w22);
and (w727, w726, w45);
or (w728, w727, w631);
and (w750, w749, w728);
and (w751, w750, w702);
or (w752, w751, w682);
and (w753, w752, w433);
or (w754, w753, w22);
and (w755, w754, w45);
or (w756, w755, w631);
not(w68, g1);
or (w760, w68, w352);
not(w23, g1);
or (w761, w760, w23);
or (w762, w761, w362);
or (w757, w352, w362);
or (w758, w757, g1);
or (w759, w758, g1);
and (w763, w762, w759);
or (w764, w756, w763);
and (w965, w964, w764);
and (w966, w965, w52);
and (w967, w966, w764);
not(w20, g5);
and (w765, w20, w764);
or (w792, w362, w765);
or (w793, w792, w352);
not(w17, g1);
or (w794, w793, w17);
and (w795, w794, w47);
and (w796, w795, w764);
or (w968, w967, w796);
and (w902, w433, w764);
and (w903, w902, w52);
and (w904, w903, w764);
or (w905, w904, w352);
or (w868, w763, w362);
or (w869, w868, w38);
or (w870, w869, w81);
or (w871, w870, w352);
or (w872, w871, w33);
or (w873, w872, w362);
and (w874, w873, w84);
or (w875, w874, w352);
or (w876, w875, w443);
or (w877, w876, w763);
or (w906, w905, w877);
or (w907, w906, w362);
and (w908, w907, w433);
or (w909, w908, w362);
and (w910, w909, w433);
and (w911, w910, w433);
and (w912, w911, w433);
or (w913, w912, w352);
or (w914, w913, w362);
or (w915, w914, w27);
or (w916, w915, g2);
or (w917, w916, g2);
or (w918, w917, g2);
or (w919, w918, g2);
and (w920, w919, w76);
and (w878, w433, w764);
and (w879, w878, w52);
and (w880, w879, w764);
or (w881, w880, w352);
or (w882, w881, w877);
or (w883, w882, w362);
and (w884, w883, w433);
or (w885, w884, w362);
and (w886, w885, w433);
and (w887, w886, w433);
and (w888, w887, w433);
or (w889, w888, w80);
or (w890, w889, w352);
or (w891, w890, w29);
or (w892, w891, w24);
or (w893, w892, w362);
and (w894, w893, w69);
or (w895, w894, g6);
or (w896, w895, g6);
or (w897, w896, w352);
or (w844, w352, w456);
or (w845, w844, w763);
or (w846, w845, w58);
or (w847, w846, w80);
or (w848, w847, w352);
or (w849, w848, w24);
or (w850, w849, w362);
and (w851, w850, w71);
or (w852, w851, w60);
and (w843, w433, w73);
and (w853, w852, w843);
or (w854, w853, w362);
and (w855, w854, w433);
and (w856, w855, w433);
and (w857, w856, w764);
or (w858, w857, w19);
and (w859, w858, w764);
and (w860, w859, w52);
and (w861, w860, w764);
or (w832, w796, w456);
or (w833, w832, w763);
or (w834, w833, w58);
or (w835, w834, w10);
or (w836, w835, w80);
or (w837, w836, w352);
or (w838, w837, w24);
or (w839, w838, w362);
and (w840, w839, w71);
or (w841, w840, w60);
or (w820, w352, w456);
or (w821, w820, w763);
or (w822, w821, w362);
or (w823, w822, w352);
or (w824, w823, w362);
or (w825, w824, g2);
or (w826, w825, g2);
and (w827, w826, w73);
or (w828, w827, g6);
or (w829, w828, g6);
or (w830, w829, g7);
or (w831, w830, g7);
and (w842, w841, w831);
or (w862, w861, w842);
and (w863, w862, w433);
and (w864, w863, w433);
and (w865, w864, w433);
and (w866, w865, w433);
or (w797, w362, w352);
or (w798, w797, w19);
and (w799, w798, w764);
and (w800, w799, w52);
and (w801, w800, w764);
or (w802, w801, w796);
or (w803, w802, w443);
or (w804, w803, w763);
or (w805, w804, w58);
or (w806, w805, w10);
or (w807, w806, w80);
or (w808, w807, w352);
or (w809, w808, w24);
or (w810, w809, w362);
and (w811, w810, w71);
or (w812, w811, w60);
and (w766, w433, w764);
and (w767, w766, w52);
and (w768, w767, w764);
or (w769, w768, w352);
and (w770, w769, w433);
or (w771, w770, w443);
or (w772, w771, w763);
or (w773, w772, w362);
and (w774, w773, w433);
or (w775, w774, w352);
or (w776, w775, w362);
or (w777, w776, g2);
or (w778, w777, g2);
and (w779, w778, w73);
or (w780, w779, g6);
or (w781, w780, g6);
and (w782, w781, w433);
or (w783, w782, w352);
and (w784, w783, w433);
or (w785, w784, w84);
or (w786, w785, w362);
or (w787, w786, w352);
or (w788, w787, w104);
or (w789, w788, g7);
or (w790, w789, g7);
or (w791, w790, g7);
and (w813, w812, w791);
or (w814, w813, w352);
or (w815, w814, w84);
or (w816, w815, w362);
or (w817, w816, w352);
or (w818, w817, w104);
or (w819, w818, g7);
and (w867, w866, w819);
or (w898, w897, w867);
or (w899, w898, g7);
or (w900, w899, g7);
or (w901, w900, g7);
and (w921, w920, w901);
or (w922, w921, w352);
or (w923, w922, w867);
or (w924, w923, g7);
or (w925, w924, g7);
or (w926, w925, g7);
and (w1036, w433, w926);
and (w1037, w1036, w433);
and (w1038, w1037, w433);
and (w1039, w1038, w764);
and (w1040, w1039, w52);
and (w1041, w1040, w764);
or (w1042, w1041, w352);
or (w1043, w1042, w362);
or (w1044, w1043, g3);
or (w1045, w1044, g3);
or (w1046, w968, w55);
and (w1047, w1046, w926);
or (w1048, w1047, w16);
and (w1049, w1048, w926);
and (w1050, w1049, w1045);
or (w1013, w763, g6);
or (w1014, w1013, w352);
or (w1015, w1014, w362);
or (w1016, w1015, w104);
or (w969, w763, w362);
or (w970, w969, w352);
or (w971, w970, w362);
or (w972, w971, w352);
or (w973, w972, w362);
or (w974, w973, w352);
or (w975, w974, w36);
and (w976, w975, w926);
or (w977, w976, g3);
or (w978, w977, g3);
or (w979, w978, g3);
or (w980, w979, g3);
and (w927, w83, w926);
or (w981, w980, w927);
and (w982, w981, w55);
and (w983, w982, w926);
or (w984, w983, w407);
or (w985, w984, w763);
and (w986, w985, w926);
or (w987, w986, w968);
or (w988, w987, w58);
or (w989, w988, w10);
or (w990, w989, w80);
or (w991, w990, w352);
or (w992, w991, w24);
or (w993, w992, w362);
and (w994, w993, w71);
or (w995, w994, w60);
or (w932, w763, g6);
or (w933, w932, w362);
or (w934, w933, w352);
or (w935, w934, w362);
or (w936, w935, w352);
or (w937, w936, w36);
and (w938, w937, w926);
or (w939, w938, g3);
or (w940, w939, g3);
or (w941, w940, g3);
or (w942, w941, g3);
or (w943, w942, w927);
and (w944, w943, w55);
and (w945, w944, w926);
or (w946, w945, w407);
or (w947, w946, w763);
and (w948, w947, w926);
or (w949, w948, w352);
or (w950, w949, w52);
and (w951, w950, w764);
and (w928, w654, w926);
and (w929, w928, w433);
and (w930, w929, w433);
and (w931, w930, w764);
and (w952, w951, w931);
or (w953, w952, w362);
or (w954, w953, w352);
or (w955, w954, w362);
or (w956, w955, w61);
or (w957, w956, w13);
or (w958, w957, g2);
or (w959, w958, g2);
and (w960, w959, w73);
or (w961, w960, g6);
or (w962, w961, w94);
and (w996, w995, w962);
or (w997, w996, w94);
or (w1017, w1016, w997);
or (w1018, w1017, w41);
and (w1019, w1018, w926);
or (w1020, w1019, w55);
and (w1021, w1020, w926);
or (w1022, w1021, w79);
and (w1023, w1022, w926);
or (w1024, w1023, w81);
or (w1025, w1024, w352);
or (w1026, w1025, w33);
or (w1027, w1026, w362);
or (w998, w763, w362);
or (w999, w998, w352);
or (w1000, w999, w352);
or (w1001, w1000, w362);
or (w1002, w1001, w352);
or (w1003, w1002, w997);
or (w1004, w1003, w927);
or (w1005, w1004, w362);
or (w1006, w1005, w36);
and (w1007, w1006, w926);
or (w1008, w1007, g3);
or (w1009, w1008, g3);
or (w1010, w1009, g3);
or (w1011, w1010, g3);
or (w1012, w1011, g3);
and (w1028, w1027, w1012);
or (w1029, w1028, w80);
or (w1030, w1029, w352);
or (w1031, w1030, w29);
or (w1032, w1031, w24);
or (w1033, w1032, w362);
and (w1034, w1033, w69);
or (w1035, w1034, w997);
or (w1051, w1050, w1035);
and (w1052, w1051, w433);
and (w1053, w1052, w433);
or (w1054, w1053, w59);
or (w1055, w1054, w11);
and (w1056, w1055, w69);
or (w1057, w1056, w997);
or (w1058, w1057, g6);
or (w1059, w1058, g6);
and (w1062, w76, w1059);
or (w1063, w1062, w997);
and (w1067, g2, w1063);
or (w1073, w1067, w352);
and (w1065, g2, w1063);
or (w1072, w1065, w362);
or (w1076, w1073, w1072);
or (w1078, w763, w1076);
or (w1079, w1078, w362);
or (w1080, w1079, w352);
or (w1081, w1080, w352);
or (w1082, w1081, w362);
or (w1083, w1082, w104);
or (w1084, w1083, w997);
or (w1085, w1084, w41);
and (w1086, w1085, w926);
or (w1087, w1086, w55);
and (w1088, w1087, w926);
or (w1089, w1088, w79);
and (w1090, w1089, w926);
or (w1091, w1090, w81);
or (w1092, w1091, w352);
or (w1093, w1092, w33);
or (w1094, w1093, w362);
and (w1095, w1094, w1012);
or (w1096, w1095, w1076);
and (w1068, w27, w1063);
and (w1069, w1068, w1059);
or (w1097, w1096, w1069);
or (w1098, w1045, w1097);
and (w1071, w1063, w1059);
and (w1099, w1098, w1071);
and (w1100, w1099, w1063);
and (w1070, w1063, w1059);
and (w1101, w1100, w1070);
and (w1075, w1063, w433);
and (w1074, w1063, w433);
and (w1077, w1075, w1074);
and (w1102, w1101, w1077);
and (w1064, g2, w1063);
or (w1103, w1102, w1064);
and (w1066, g2, w1063);
or (w1104, w1103, w1066);
and (w1107, w55, w1104);
and (w1108, w1107, w926);
and (w1061, w60, w1059);
or (w1110, w1108, w1061);
or (w1112, w968, w1110);
or (w1113, w1112, w1097);
and (w1105, w16, w1104);
and (w1106, w1105, w926);
and (w1060, w12, w1059);
or (w1109, w1106, w1060);
or (w1114, w1113, w1109);
or (w1111, w1108, w1061);
or (w1115, w1114, w1111);
endmodule